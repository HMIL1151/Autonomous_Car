PK   $xXkU���  ��    cirkitFile.json�]k��8��+��Y��I=��t�,6��t����PzP]�8v���c���%%�b�T�{��.6ݨ�,�������"?��;�+��A�����V7,^���C�<�4\�6��/~?����O�����A�A�M�Wu�4-CUIEeD9�,��@ĩh�2L�$)�"\�ܾY/G`d��`dT���dT��dT�����a�9P�"!s�"�EJ�@E��́�9�A�(z�$C(�PI���,��=\�!z�$C(���A|��o�;�;��2Ƴ4�D��`Y��a�iڔ)��`\u�����b�����n�dq%,`B� jB�U���2�e����K�yz�'C(ل�ʤJE]�@��R �%�uP�7y�4�j�A�z7���D��8�8��� � �!��wOd�0��wO��=�!z�D�P,��B��� �����։7�Rn �� ���.&���t���M�GԸ:�-9�N�0b�#Ç�{y�f�<AU<��as��*G.H���߉pˎa٩�vk;(;�e��sX�q����]X���vPv�.,"��"����]X�X��X�A�1,��H��K����cXva�bm�bmeǰ��"��.��ʎaمE��]���ò�/t��cpf�������(����:� ��`0p��������?���Y���/.��gX~�O�r��m`�10?��l?pƁ�����Kc���Y��ӯ���gX~�O�m��}`�10?��<��?����^k �8���c`~z��~�7�W������?����^��8���c`~zM�~��ˏ����@`���,?�#���?����^�8���c`~zM�~��ˏ��o����]���Zg��yFi�S�=��.��RZ/��Z��<�5g�eD<+�L�m U�,qInl��Y}��{f����ǋ�gV'�n�|yf������KwgV�͘Y}�/c��Pݎ�w�^�����g��[��{��|�ޤ����g��w��gli�[���6�����glݘ[���ƅ����ǉ�'��'��'�/����Ĵ�9n�4Xv�YKl=�0:�����\!�NNH���n��uZ��m�%��Kќ��-�RZO�����>w���O���t���a��|�"�P���a��0�@@�����0uJAF �N7�ԩa��:M!#P�0�a���@!�qa�,p��ze"'X�f���B�U�@�:��p�pR���ᬋ�"��9��8�����<j[��{$��UE���(�^��	�9,���zA'X�8�B��~V?��:b5�,��.�f<��X��	�y}�4���)C�����aդ����51+ϑ�246���h��(�Ք����ꃫ�[���x�4hW\MM�ƫ��@���j��`,0^mG��WSc��*l8*Ю>��:9�Wg�Q�v������X`�j�
���������pT�]}p5�w0���ꃫ����I���O�六E�������O�e���a����zyak����"m�'����"��E��O
慭E*����4�[��i[?����!<,Ҷ~�1/l-�CxX�m��d^�Z���H��I˼����a�o��e^�Z$��H���˼����a����J�O^fH�a�����yak�I��"m�'/���"���E��O^慭E^	������[��i[?y��Y&<,Ҷ~�2/l-�MxX�m��eNl��9P�}��|y%����2I����厞���� eb��|$ ��j���H ������ (���%P&��,�NB�`�wj��A%Ɓ�v�-PYB�`|xjS��%D��x��n�zL�Om�Y ҄��x�����M����P�����E/vU|�8����l{��+)�,���+"����W6����P�n�/掼��A�=t���� ��T�$@ h'O�r{�o�  � �0�@F �^ �� A��z #P/ a�� �@@� �� �0@���ڸ����QH� �,v3X�F!@N���`�4 a8�b8�q�  �����QH� �n�����8��q�  �����QH� �,�sXG!@N�8�aq|
	  �F� P-@hTW� hW\-@+�Ѩ@���j �X�X=�F��W� ���a4*Ю>�Z� 0V�Q�v���" ���b�
��� ����hT�]}p� A,`�F��ꃫE bc�0hW\-@����˔������\^����H�zJ���]��i[?���6 8,Ҷ~�//lm@pX�m��`^����H��Iü��	 �a�����yak ��"m�'���& �E��OJ慭M ������[� �f�O^慭M ������[� i[O����e��i[?y��6 8,Ҷ~�2/lm@pX�m��e^����H���˼��	 �a�����yak ��"m�'/���& �E��O^��v� eb-� :��z�@Ϣ8 �Q^��� �E�: �Q&V|/ ��L��^  DG�X��D  ��ީ-vK� 0��{�D  ���MYK� Q��S��� `0^<��g�  ��S�[� `0^,0^,0^,@C	�����Y ���0�v ��`�8����(/:�� �Š�, ���Z��é������4V7��W�7y,�e-�b�+��FV7������m�oEă$�"�m�p�a�V�d"O�Z��ެ�7�(MsR�jOnM3Rӂ�tHj:"4�O�,b�F!o��e�r�8�Z�AɸlX��q�H^�Z�8٤{;��Oډ�d�N�)Z��)MO(��5Ms���4��f95M�'j ?Ѵ�(��E�)��Cb��e�(��k���wl�Ӿ��������J��9�OF���E*2�@�H�i]���E��>}��u��uj,�8?ѻ/��߷�Y��By��)�.i}�܇�o�cV�)�8Β�A{X��ʽS{���:5�O�q�3u�8���D�A�ݿ�MQ�ۤѭ���f����I�Ht�y$:�t�qV�Y�br�N�8��,�o2�D7uƉ΀:�Dg@��3�NCu���`}K$@���&��L�����D2�̀<4"��̀����̀�m�? ������������M��ķ�*����K���"Ҭ�K���ޑ���eyǤ�1ϖ,{q�0Y����-�b����i��)~����9W2	�+6@ئ�^ְ��_�,Ae��b<�]_ �,A}
����'B�D89�s�2��0���'}�q "1$�_ @GN �,A!a�^44ZN"uI~���	:	�
:	�R
�a�mE���t��t�e��J�y����~�}���C�7��F���MdA���&� C��sY�!�#��,��1�Dd���m"2D�6��?b�Ȃ��MdA��Ҧ�-D�D�O@�d� J��ɦ� �P�t��8l*���i�j�1bE��bSi"m��2�5���p"6� �v�[#M��aSo�I��S B3c8���9 4�1�Ӯ�< ��B3c8�z���`�����h�DZ���-��4!Ŭ��IK����6!��( p�u��U0Ix�3�qx ~�s�qx�a�YN�&ޯ!��Ã���rz5�~�{�~X~�S���k��� ���FM�_C�������i���8<����,�K�����A��g9E�x���<b?,?�i���5��qx�a�YN���w�	�y�2uċNA�m�>16��!�<�<1��!:3����������kbl�NI�m�216D�%`��󗁀�S0C�9�@@���	���<e  Ɔ���vn2cCt�fh;���F�)`��s�����0C�y�@@��L�y�yR0cCt�fh;���!:O3��S�������#bl��S�m�16D�)`��󅁀��0C�9�@@��y�g�<�{������͖�y~��l���Wϖx����i��*�����3��zg֧��XE;����uf}c]���������u�s���T4������[g. ��ͭ+s��h�0����h@�Ds��\ �'��
�P=�\�?�ꉜꉂꉂꉂ�-S=QP=Q<�ΧJ����M�2;����.�����И-�����ي)��i��]� 8�;��P�q>�w7���x�o���Zo�hx�2 .i���v��A�����3uV._E{��J�=�����ޡ��y�%�.�tY�3]���^'��t�k�[��Ξ��5:%�N�S��䘄�!t���5��!��+�o��[Қ+��e�Q��2;y��P��4n���fP��(8_fy��q3�x3D)<JL3o&�p�ov��9�A �8i��2�}����HO �8!��g	��ƙ�!�Inf_O �8����Ⱦvd'��Tl�Jnu6����M����ht���y���y).E�x����pI����Rb^J�K�y).e�|����k�(���mqf�ͮ����lڲ:l�Pѱ��(Tϲ�q�j֦U��!/Q�����Qle{҃�g(�/5�ױ���B��$+ �����<�
�S�����AN����8�����T���Bpeqo�u*�k�y�Q��D
W��FXDq2���$��*����s�m#�������5�Wj�|*wu�4f^����B){���)ԛC����2�^���oַ,���~��n�~!���[k�����������oŮ�5W�g�����N����JO���wu���]_]�ޕ�G��_���
��r�����~����O
wuӖۣT����温��鳃���� �yO�C�s~[�۲>=����΋�1�L.].P&�?�:����O�s�+K^�����@�Q��/�A�7!k�,����sl�sN����,���9�h�r����ԕd�N4YGL�a�u©:���Åt�F<�H4U��k�'^�*_����q:|�҉6�_/]HL<����Ù(h>���棛(h>ɉ��5
�����Э�L�3�Z���rg��3]�V��Hvrar����1��˙S9���x�r6�ؑ�Q�.4:�ǱX��m#�Ow]�p���[�!O���j}��4�'jh�򶔁����Y�e���oԲ,��FFmW^~x��Uo�立�W}ݸ<l�8��7j�U�A6Q�Ta�dU�q_W�V/me&�*X׹
�Q��L�����de܄�?�{�{x<�UΒR��:hҤң�T�2"5ʈx^f���M��W����ge��/��;��~�mΐ�I2�3�)	5���6ȳ���d�I5��.L�Sy8�O�<��J��8�L���V1-K���+YՉYP~����k
5�mZu��en�#�����&��p���P����Y}6(�������j�!ޔ�7�r��j����79��z8��i�x�}^�u��u��J�w]o���2�x�HVA�#=�L3�%��*�8�q���z���VDe�iR�G,�P:�M��U��n�<,j���y�a���w�j��l)㼬E͹H'=,n�,	+�0֖W���*�(�*mU��{X��z�z��4WGyz|�ӿ\}���]]���W������C�J������:������ܨ�����_�v���-7;�A>��$���s����r+�S�3��k5����������.S��]~�zC�����M�7��W��Q�QwLǺ�g"�Xu�:��$̆��|�6�E�F�"��ϸ,�4U!#)KcS��vF;M�����F'��:It���TwT���˒��yx��l��o�0k�E�c*�#���L�g㶉�:Q)���:I`<P)x\�Q�����LN/5�fz|0��u��I?����/b4�J��p>�JO�W�F�_z:�ˏGOv�wM��=핗�2�pyؽ����U�������o�ӽ~j��<�~t/7��뒩q���d�ø��sp�����e���\��<�>�������KG=��I�^Չt�����H]�S�pz��!�����v�n�P���Ez��
��36G_��������N���}��z�������}�/��ѣ���V�첺���"J��cv]b���tA����bi�K2{�I�]���b_c�e��L�R��g5�R���Ck`WNp�zt�PW����G3�W]��k�T��♏�%�T�k�ё���x����ګ�9��\��7 Gń��Djs<&��bnn�����<v�<s�y3��t;����e�,��|��Z��3��U��L3b�3W�3��E� [�/�ɱ��S�<�����Jd��E��9.8q�}b���>Q8��b"��X��/�pk�/zT�RS�.I]�b����*tPqN,<���b�3���e1aOB�(2:�J�եx|��N���_P�щyXG56�u����[v�m�ݝؙ�L'f.�rY(�'z�dI1����*y�y�v� 0��*�U� p*�\x@d�ϖ�Ƌ�"�������[��i�a�ia���q��)�Q2�X�5��[�X�?��h.+�=���.�r��-���&]�XR��Y2e���%�9K��YR����b�Ko5*�F��bs��/�nŸ�ht䡎�;ɐ51+�I&p|�sw�L�3W��|"�%���xj�nŦb�^M��ni.O�)�Z�Iyϱ�e�߲���=���o_��[� �������PK   $xXo�>��q  �q  /   images/2cd737db-51bc-41eb-8762-f3273c40eae5.png =@¿�PNG

   IHDR   d   �   J���   	pHYs  �X  �X{�M   tEXtSoftware ezgif.com�óX   5tEXtComment Converted with ezgif.com SVG to PNG converter,)�#  qIDATx���d�u�+wuu���9�LO�   $ DҴ��l�Ғ�//�����o˖,��%�f	H�� #@�<��9��t��s.�}^������*LWx�{O>��+�/�xF�`�5Ci��� ��ɂpE����0�(M� ~>�ؼ�Ϡ��E�h�slyh�lz�k�.����ޏa~?.�7*f$c躴W���8��F����kX'L�{�������������;��|O�ԏ�G��Iy�7�r��f�l�)��ϔ��_��R��zmU���˶ғgsy��YX�&ē�Af\|�j��,������XC�����B����c����
�k߅��,�๸zb$?wD|roS�r�$��%����׭�u���fHL��e>��0�w����q�W'3�����/��'�A�s&)+c1fL�0�y�����xP1�O�^j���-�^�^�1C�ɰ�q���K�pq�mȘ��r�H�z�Ɉ�3��e�:��U/��_R�|U�J��g?ٿT/a�}��=�^�׻�U��;��ں��>����Q8Jl�%���3����9�}`4
�JSN��蜼a&���~���� �qj5Rg𚚘�"dN���T���yo�x@�K�m��~u�fܱ��F�շ��jZj2��.M}�W̐{|���O�aځ��]?����m���w��+������돖s$f�݊P]����=����A�g䷅�Иn/1���V�O��߁�����͙MbN'(ok]g�V!.��%�7���PO99vje��M娭.��T&��&����1_XM��T&�Z�u7��²����Ȍ<��;]�/�^��_��n���y[gF��~��a��g�`�u,�!$��8��b��� �V3b���J�*��ho��4�W��^Ĥ'R ���4�Z�X�U�V�nW9��¸��]�82�dL��Ɂ2G	l6�.�z�Q��.��'W���D0���w�_B���������m��� oc�$�}B'�{��[�j��>���7�N����oe{�!(ťQ��/m�+a�P8_(
���:~9�O����5ÙV�հ�5msAL��KHnv�Q��t�l�� ��UR��1��.�t�Ӭt��V��`8F{U%&� CA_�41,c�g���/�h��"�X��AӮ���E���A%��"�_S>�&u8���ΐ{�k�z�q���i�����-�f�ɑIܮd�_�qkj]��d����"FYi)�������I��9,-�J�8�N�J&10�E8�+��E�(ä���9�X�xnIf�[�a�K����+aK�`���]�h/c:C��L[ZfDf|S�6/�.�������'S��T��<"Ay�����>̏#�b^¼���7C�PL##����`�8�ל�L)�a��d�d��yJV9�������p����_������H0Z�����[�������Zh4/�x�������TF�\r��p�e��lƺ:7�?�+�I=�'��=WE4����ai)�^�xj��e��D2�٫a��ӞP�?>'
��M,a8��A�#�Jǐ�]��8����A�uU��K����ك!�?�(�[��,8�+��8�N��[���Ħ�e�+�2��,��U�eQ�>y�,�͍5x��E�è0����@�W���U.~|c���*�Q���:�M�R^���"C2�)dm�I`6�5Q8��=~�vZ�J�a��#�?�}.4��3i��
Z� ��hi־>Z�E�9�ECi���9�F�/d�k!Ys1�a(� �l�P�L��T\-5�ƹ(��4*��̱83�3?���4e��$�:sB&�@ځ��2�sFe�L��,N�"ڮ�Z�I�.���nRք��8�a��	dсH%����Vem��]�z��M81<Y�3�$���i~���	���xlp>eyݿ���	*��u@�o-��S�#�P����U����ؤO�0���2Md�PVQU}7��~ e�b��Rq\<�.�~S��ȴs�V��*$��]��OO]Ƒ�qaC�5e�p�,�V�,�A3}�@>.ǂ�妭��ýsT�0S���3^�8�������Ճ7.�''/#O�t�.���!l�p#�l�[Mv-ҞLFP���>��z�S+�S�Ȑ�Qgv��(�6�:@���ذ�$�a\�tX�y��'����E�ꮀ�j��3.���|D�������[�aH����7:E� =�DzQ_��1b�9�ڱ�DF�X�8^�Ua��nU�e�HT_ ��U,c^�����(�����dZ9�a�[6���5X��~d2i���V�l��]"�↨�Dj��S�+�4�n�����_�4��f����m];p��	�	t�&#qE����كjFT�m����;wh��xbY��E��*Q_��\ex�^�>7�ya��S�6�`]W��w8J�?��/�]�82��2a��F	J���e���g�+��p5v�� d�zQ�әt��h�%�ؾ]�ӈP(�hTcHYY�_�hjߊ����zTK3����VR.�������.�(�b2��J��s�$��(�?��4�܍߹k��c��b������D�j��� ���h�C1�4Ӑ��(u�p$�Q�ʫܕ�(��Qj[V�y�Qf�b���Q�j���)T��g��t�θ���lu�ԘS�ȋJ0>�*�/.Y�7��ۡ��P�IV��h�L�+/E��G=�~�6��7�T�dX�7�Ջ,�3�7S�E�dõ05x��� >��M�EgS޹2�hքx&��o�����3�΀w!��t^���"��b|��G�P]ی��!�I�ӱX�hѼ�����_oǀ�����:3�ş������_|�nL�cP4-1��x��t2#J��,�d`��sIu�O���Y����2â�-��T0U�`^Q�~������?��K$k��2m�{��a�N7***�����0����d�R�f[���K��8~��X��.Tմ�>?.����e9��@M��><0����(�a������>�?P�Դ�U����R�5)�8}ދP$�&�҄��sJ6�d�(�:'�;�Y"J�_��:0��s�BPD}\Mʛ��ٿ��s�S��B�������h]w;*�u��o�^�Ao��Nq9�1r��I�<8{��ܝD<�DU\}G?$'�/}�&W9��=7(k"%v�����	���,�a�-�9J]��o�5s��S�B|#Ô�+�n�¿Ӵ�Nxb3��i�N���X<m ��/���_�f�_��d���2�_SVz���jS>�7��x83
�i8�er��X�#��I�Y9���4>@�/��0eՏ�,�h��\�_w�6��K���G�����sd����Y���T�[݁���3*O�xLZ)�ц������w�@\��i왨[����ʴ���B	��(5*�9Yۅ�����e�,t
9	��4�9)98��%��d����-x��i7FR�c���|{0ZQ�O�%��y^�d�Z��YA �U�m��o2%�H8Eg���=��Wˋ���-jA�F&٠��dm�|ҫ��Z+�rt��&��{�*%��)�t�?�s3j��sT�����R\q��.%Jq�P��;�2�GQdY+Sf,�1+�������VL��$�v����o߉py���rL�i�J����������[�8��r��|d�|�����&�n[638RjE|F����~�,���\/���%��>����)�rb!N&�^h����>Ҹa���>�jʚ�E��u�ߜ�~w3t�)6�s��
;��nI�&k�B+�[���s;�x��E�$G��\�tg�E�9�Xd�p�k�7�9�:sR�7c�xƦ���C9Y�<t�L��R��4�(TY�m�d�ErzlJnX����vqE�ߧM�¤��_
�CjcU��?��)�Z��F���9e8��I&����7"�Ί��O�4d���$�6%�ϔ����	�OŲ����+&q�ÏjG�� �Xg�6�$� OZ;�<V�0�̐��Ϣ���6��z�A˖�sX��\������|u�]��_��0'���qiZ��8��'��cq�"�L�T�����PT�}�����1�D-��XY�WN2N�jK���FG��r�:�co�/�k$<��MQ��ϸFqWMk�<��n1{#!�N����~|�ӆ��*rw[=�{�,.M������X��;�� �~�y�zK������oܲ����F����qyҏW����Y&��@����{v������僸��N��85�A��&"1��}�o�/���fū��3.{�V�����\3��V���h���^u��@5�4~��[��v�GQQ�CBJw�{������h�C��]� nq&��/���	���i��۾�D��79�暑)b~d�ZY��~�����=r'��{=~��ױ�wX�m�b8o��R~_�syXf�ya?��7I�W���1���{qcg~���xJ�<�$*����AyΕ�-��/Wҗn؈�/���=nSף�Ģ���ٖ3��W׿��Yy�!���,E�����:�АQ�����f�28��V�d�[8��p�)J��y��$ �ު��CD"��f�Z�vW���Vly
���Z%F1�XC1u��v�W8�~����~���Ͻ�?�м�U�A��P^b������$s	�e���G���W�ƍj�S�Xc�I�RE�l����-Aյ�9vQ�X_
+q�xۋg����Ŕ 6f���5�5�J��+��ɘOo_��)�w�����0Z�|%%�������(--�PJ{�lۋ��!�1$g\�4�*�E1f���uO���Ҳ*T��(3*���+��y�6T)낡���hQ~2O��H�s�"���f5��ֹ%>ƙ��ۋ_�Y+����n���*�'<���5�2591(.�&X�����~�
����qD����FYi7�5���ʛ���j����|�<K���	��*�98Ԕ/U�iH�&�Zy4�L��V�(#*'�[��i&��Ab��E��ň�AQ'��VM����h0*L�\׽f*�?���N1��Мd_��D�~����R>��5�Z-����~"q�,�����*��G�Y��W	�=ј�r��o\]ĕ�����#%�ۧ�j����\������Nq�;�+�k�^;x!��<b� ���w��FD�w���j��!�SJ!�S��&���p�\r��b�0r�8��F���p �̿P�Œ�}]��'�L�;�O�O^: E��2���s*��s��)3����3�"��R���aa�o=��X2�� !#�X陚r;B�c��ӭUZg��/J���~�������ij6]ۂK!~Ef߽�M�	���iF����i=ʕ�ŕ����F�O�r�!<(����F���Sr��Oѽ�>�W��g�TO�����x5� "��`�(k�ܸkj\��{��o�(�$z��#�����"���	qEP��z���^%�cx�L!�c�siǘ�SǑ���Z3��Fÿ�c��C��߾ye����ڎ�^�>�<:�߆R��2��q��k8?>�wc������?c��<���H�qT�[`4[�c�7��kq:^��!j�ݥV{?���I�|�
�y�mE���H��6J���P_%��R�E��ӣ^�I��uI����iҲ)��7u4���J�E��9�X��Z�TsL�����E�N�@V%�I��}�d���^�Ӝ=��(.����Yh?O�=��d	�z�[��'�%�8�<���6Yzz�KKG�2�ej%����Ĳ�P���A�S'���ރ?{�Z}�/n݊�z��]��XU���l�§w����]|lC��q>ea���rO_T&/E�s�{���|nZm\!��1X|'�Do��BAԍ���K9]�ɚfĸf8	���(oG�xnM�C�dM>R|G��4?���Qu#&���o]�v�Pщc ��{{ڕ?��ev�I�$Q��k�'��`��W^;$���߾s��MW��c��i7���tʹ�J-5;�8�k��eD%�0A�8��R p����o��]��z���ӆ���W�ʭĘ[�K'�֮&1>�R��M�P��s�����Y�WOH9�sA7z*�7�7����S����,~A9t�Q"�̸A���UI��Jaڔ����٩^|�|/+����m�老C�4��k���"�K6�:��p�iW��\�N�0���C9��h4gR��aNTR�OVc𬴰H\z���Qlo�뉦0���p���X\|!��_}�Q1|S1�޴	�����ӧ��W�Пb��B���t�)����z��t�*��2٣9��8Y<h�=�[4ZSb���F���/����h`�ɋg�Dw��Dx�| ������и��ƊM2�0]���0=� ������_�}5E''��G��C$�������防×��rv�����CI���58�(�_��w��>�DG�&Եl��dE�;���c2�L4%�󚼤���^F8��)�z� ���&��"����B�]��7���C�B��T��E5{��
e�"U�_�|�I��k�Veб�V��:����]Ės��Do��f��dF�-�O�&�u����=���XQ�Z�6m���'0��⥐V�M��*&�8X�z-g!e1����eI�?�m�]��[׈N�2])}Zd��cJ�3,O���k59�3�&#����5����7���/���^aƎۿ���v�DZ�������a0e�ج{����^�6u�m͍�E�H$��Q�����tm�7���ވ1�@��fl�D,��w��J�+���l��z�2��wN������)�͕I��*�m����������X[�߭�"�=(1FCQԖ;��c���þs�U�C��P�����TJ����醵X۽M��4.'����R�4Xp�vZ��bkV0:epV���nB�)���8hgl^)���Pj���ޡ���,:���[E$/r��Y��>���������Z����YPJ������|��볜��o�$� ��{q��p[������ee9Y%��c�*��
K�%�󘲜��l�PԠ�ݥ%�፼��UWUʿ��*yA1�Wv�Fc�	Ix�p�����7��VL������(���>"����S�L\񅋹�tZ3|�[��Y/��˹�C�tG�vx�.�}������`�
&F.a2�G0kE��{]+�V���a�����lZL��3n�\8�r�ҙ�bJ��Ă��،o+S���ݿN5Y�"a�N:$�&2�7ٰ
���}cH�,�eL:���u"����զ@C�n�	fd�Ǫ�{�N��������^�V�����*�W���ɬ��Š��Mba\�R�3�N�����7 !��:�^R������bV��ad�^J�+�`m�m�P/W>��6x��Mh�ڦĔ�M�Us��>�]T�i�Y�`*����ѳo!���~�t�����C����*1.-ګ�9�yCb����c8�����ء�'���)�c8E�3LQ��h����<?���=�L3;y��V�0�!�vI�O���L\Fe��0蹂��^<�U�����qb"cŭ�Q4�	��i3�\�9��.^�=e9+Mh�9�"�!�U�j�����տ7����\��l�t��X8��0j͞�ՋY�+rU}�.k8e���f)/]4���E��O(��:�� 8;g(WC�_ж���c��C'�F*q(Z�cN�x,7U�=}�	��?`�]�ȟ]��YJ����\�!�+��=��4��X��w���R�%#܎Y%�T���EKQhCX���O��i��.��u�Y�x_ؽAV
����B\����C/��T� 4O���h�Ӝ�N{ m��0�E���.�J�ˌ�	�3��+qE9B�T68�㯝x_��}��-����Eh���G�Lɂ�^�<�BWU%j6�d�"�����i�����n�p�Gz�j��� ��w0��8ӥ�E��sm�m�bE�g�g���I_�KKB1UeNĶ���a�'�W�Њ�Ez��v��+n�U����ӽ�pWJuű�	iN1���1Nhf
!�E� <ӏ�ou,^��� !�i6�5o��H(?�v�B{�^:t5�(�*϶��|[�!y�#b��Sk[i��'�i��б�&ɏPtf3�9�&L���_��I�ŗ0�:c�Ç��jl����؈HD�bd�Yk�n���=�3�r����Şz�rGs��CҴ�8o��������-�MR���֊���d�bc���6�uXR�"���K2��'r��,b����]�ޟ�K%�Y8A��o�;��3�;)3�=���n߈Dx������`$�eh�؂�u7�F�P���T�;D���OC���K��˥�A]�͂��0���Ӳ�J$a�|�� O��f�U �6d
���2��ě������]�]���|�Y�׭�4��C�&�mz��rg�nu�C�c��vIg������qɂ�r���Ȓ�<�9��]�B��`�=��$�&)l��BQϝȸ�VU!�bN%u��*ڱ���^ZC�K�B׮}��pZިt�1�n��5ɰ(�b�7o�,���К?Y*�r�\Y!�&�����7%��X��C�*"�-���C��ݒCg��rǽ��$�2@�bQ6�t�XGt(�}����,��)�3ׯG�R��!TF��RY��i�k�����_gBk@ �Ƽ�@��z�ח�"�P��� �A0�A$G�g�ZC8;�Q�����d� ����a�e0,�(T��7P%f�d�:�d�1rJひy9�2>�OO�j�35I�g�߫VL���@q�ʹ~I�2�lf�~8��׹E���\JWcؖA���6�D���S�b�(	�@]�"j�N[��;�o�,<��1<wb��E��AS�z��:�^\؋S�2��b��h���	�̿|�&��Tc���A,=����<j��H�ܪV_D�����B������!E�>��-x��9��bI�r*\8(J�r��i��+�qbԏP2+zc4�P�c ���}�e2�u�RY�FI��Ա=�R��狪kJW�ҝ��'����cM�w�N'*�|E�׺n�,q:�"v
�ѡ��?��_�T>DDq�D�o�����G��D�	'1|i/����R�Uۘ{��K�����s���B2�ŗ����L��F�P��TΣ?��Иbʬ��Z��U|�y�i1��������q��f\�g� r�R<�Y����JN[�6wwng�Ą��6��O���0)E<*�n��j���ܜGu��S.�JY[g�#MF\
��S)Ԋ���\��J��E���F�m �O���&8�͢�~_ޏ�}V�T��̎���������������P�I����9��:��QD�c-��ڍW/��̌��X�L�V����9��^���������+-xl��D���lbQ�~eĀs>,9(2���wYQ���t��:[���98G��ޅ̒"P:�յ?�aC�#���
��/�)�}<~�$Ք|�=\TFC���PրoxZ���6�_R��"��������U0L��1DS*�*�u�ƜU�/ˬ�� E1e����<���mk��)e���ӂ�λ�51�t;��J�e��Q^�Mq#?��u{O��u�c� U�3rGYu�Dte�u0Y�72��k��g�6�-��$�D<P ���"cJ��`��'˟XֹX��l��
u|�7u��b<`K5��`�&q^&�w�����)	�Lfl˴`[��.�hΈp�
�h���e$��iv�a͔�e�:򕔽��Q��2��t!�b��,e(svA_�LR�$K+��4�b�����QKiC��4��D-���q,w�Vu�f{]����)�({�r��G�asNnOF����=c^|9�|���hɂ�=��dMI�bFYok������~{���옪6^���W8N�l-W>;�|+�K��2exH���C�,�Ȝ�!:��>�L�O�3�ɔN(g�F!+��2HEF\���=W��
�������sq��e-q�7�[�#��ҥV�n�u��h��ԗ9LdK����倧L��1��a����2�D�dRQ�Ux���t��b�m�W��fK�&��1�8��)�E��L��R���3B�E��{�v�b[y��*e�*���rh�c����×�������M�T��hi�(u�Eɮ`m ����OH+v�]��!��Sk:�W+�L�R�{bnN&�G  ��҂�]h/t�f7��U�Õ#�4�嬕���&p�o���+G�1�)~�=���ʱ~���j�fC,��ӯ�y���p19ϦO���B��AX�a�n�)+�
3FKQ/,=��Qq��j!�Eq��:�^T�%�G6��UE���u��s��z,�z�#�q�7[��ժl�ڀu���>>c,�C����P��7�m��h����Ƕ*#���"FUZ�r��vJ)�{���U�Ol��~�X�)��9g�G2���R=��(��zh<�����V�U���uk�N���X|����Z������-[$V��&[����#�+Gwc6����_ ������ �&���x+Z5�-Z�6��в�5��������Z���k�.Jӛ2a$��ݛ���=p�l5���Q��%��KP�&���~�f1�mW���rJG~e��a����yv{#�\-��b�k��g����=un��͛��ы���S����]Ꙕ?���+����]����8�*�*�p��eƬR�.�o4[��=��I�,�b�Ty�~�����ֶ
��3�/�Đ[:�
�ۦ�ei��C�DH�'g�X,���aͦ0�G��Z��5c"
�3�����	\cv���h���h(l�\q�E'��4��R��$:��+%reT��b�7[$�+�My��P]Qt���!_�k�����ա5�O�:�p�[�L�/!��FB@�<3�7I��:5��q<���@L���K)��I1Eo�  ��ҙ����V����Dc�g�W=�U1٬<�d������5�2�l_.����b�I���L֢a`T�q&��9�,$��Br.��d�h�ٞ1���J�psG�o�;�?�����$j:� �S/�hV�'gf�&+�c�,��ݨp*g�l���
I)�=t� �$�ZC��QȦJF7�z�VJ>EY�J�&�N{��u�64��m��14(shp�t�@ ��b���i�6�J'�U�	�T��H<������Ԭ�xl�RXJ�i	��:W?���粪s�&�^���\�S�	ß��n��/U���èm�H/1�9̬W�{H�l�\x C�R��Q�B(9�,:6���)E��B述��.��pK�Q�����XSf��_V�.���L0�+O�f�&�#��Y/ȝ-��$6��)e�D� �a��� Y��[ެ��\,��!���RDLd���x��blԤ������;�+�d;Z���O0�Ƌ�Zt��`>���N���+��{�w�U��*ڷ�,r��W��=�mV�� �.�J�Mf%�|�%���i�(X�u33��B1B4� �/�h�w���d��WYd���Bf��b���#{����DFrKβ�������I"K`�����\ȿ{�0o�6?If�t��z�g�S���JY\�����<�@���ʷr�"E�86�i��~Ά.�������Vt�chS�#��2帐l`��:+�Ӊ��q�I��`x�d�^�թ�,3���o�>aN�Ъ1E�p*�౦�u���hn^�$�q���x�~,���C���G���$HC3+��8w�/SXg���}1���66�*���8L�D�������7��6���5űYD�s�l�Q0����.'����b˼"Kj�a�K/��H��ł�CO�c�ֺ���H���z��ڗ����T���͢T��V���4�
����^�+l��0��"�0�8�79�(wYar�Z���A� W������_�,ZƐf.��c��7�U(�����3��CgD�)�I�z�V�����rnqxQ[����us<V�L�Z�v2M��2«���˩q�qD����$����^��a��t$��LY�W1���a��J�h4��#�)����<�i1�!�>ZE���Q��#=�!�:ϼ��~�J���&��X�IӮ�¡�Щ%�� lo���8�tH9>�c���R�C߆�FҀ�L�pp�_���:��<
gU�����>�9�*����`C1�S��n���g[�|�-�}�e�q�b��o�?5�g��M���[1|r[w��|.�1f'�MY-O䃛S-Ҽ�Ǉu��y�b�G����H��^<X9��5%�q�?AYy�Е��c�]H��\L�q*^>U(Ǳ��GS�:�7�G8,F%YL�ߎw`�ĳx9\�Hƨ����۔�4]��KoD$kn>Ih����[�(�0K	e�_���]j-u:މ�/;���ŭ�V��H�=��b��$Ƶ.��a�=��5�	3_H�n���ـ���1yH�QR�2�P�- ���L�(����i�W��i3�A�P"��@���!�o^\���<�Z]����%���XY��"�2����R[�%�+`�N����1I�V�)��!�҈7ϭ�~p�@1UX�rg�������)�e�]���d�3�5(��8���L�_&VڌT߳���-ܚ�Rf<�(��Z5�E[$XW���h#	����b���4�Mݹq� α��Wvo���������J�Vo�}�a��"����:)�(��+� Բ��<��XDb�RR�غ?����y��������E�X�1��(�yA����`DĐ3�����D=�Fu���rH�ɮ�)�cO{�0����J#����C����+�,W���4T��Y�a��a�a"m�h�I�7i�����MI������S�K��Bk�#����c/�{�G�|Ӏ�ә4z/���Cx=R�X� ����n!pu�]�����3��J�'6
1)�v�℀{Ԭdn��'/���LtwL�*\m���{g�b�0Q,�  N\��7#5�P���йn�˵�	�w.�}�G��n�m.��D�*�n�A-���՝�v�F16ч��������F��P�ݻ'����ː�,���g��	e�P�g��Ր���@�.�UIk�+���UD��9���x�j[o�}��,�m�,�-]MJ�W�J9���>v�m'.)�A=�G�7�~��U4'���8w��;pCď��c�26�5�Bܮ�. �
 ����h�RC���aT߮�j'/EлWF�|�_�-�.�99�(��Wߠ��.1�	~��Z�:��URB�3@��	I���Jq �!���Bk@�g�Z�p�Y�b/̴�)��_��z�J���	��Ё+���͝~�]��J��±�N![��������CP-��s�]/ K��5��e@k̎YM/ւ�W���?�KϜb�}xLT����|�g�nEC���+���#�D�u��N]�Y�1�k��J|Ɠ�$p=��ްH��ݎ��_� q��4���kd�ټ[��߸��
x�bA��1��*�⌭+��! ����g�/�ļ���Bt���dawV2J���+�|����֞��r�U��Gʡ2,�8���#���Z�
�&���tKH�
!O���G�|׋�Nl��}x�ET<�͖�ͥ�X�"�t����f��觑Җ�6� ��պ�!ZY{eǴE�+�~�su�EY���Ν�������_2�q�0��ы�������-�8�S6�Vc e�_��78��u^{S;j�7H���3�}'�/�ꊡb]!2/N���\���>L8U�?y�]T)�7n�"���hFGk���xꩧ099Y�+++�����+�����׊"
���)��a��vE�ֹ�u]Ҳ���]����V��1��Q>���u��X��n��O���k�[7����0��㭈[������Q�a
���~�$�[)�a@�+�a�QS�S�\�R%3Μ9�o|��j������OJ�;�(����$�3�?�Ww��~z����Q�ǽ����(��i�i۶�]ߍ��a,m�p�D۾�'$Oo*������w�\��_������k8s"���O\�������7!7�J������7��p�����<��s���i��� )�ߵkWaW�k_'�A�yOO��_L�Bi��݂��� ⿵�4(f0��O�oS�6�_�^|?դ��z��:���V�ph���^��Z�R�o�iJc"o�^p��޶F`5�E���W�����آ�����?ceLd���������Y�W�փ|���H��z��>�\p�3���P�V#�8:�2�5JK�P�&{����@������g�ޥ�_��}�ӛ6J(��U����B�����Z���L�0�k_�ȼ�T(
_����c����
�4��b��@���MwJ��<+���Z�;4�.��_Af�-2�,�8g�`��}��0k�)�x��#<��GrR��DN�ʏ̤�cu-4�VV�Gd�eMUUUappp�UB��쿦��X��i	V+r����2�|!B��`E m���E�7��ꢕ��{�Tߍ��3�58��ح��{� ���V&������� .���G�l�b4dQ�,+�I؋���s�ќIg�}���Ʊ�v]�O_酻�_����eE�=���۽�J����!8iA����k���'j\k�Q�W����GM"-�˕�w�(��`��x�b���D)��a:�"�1%���hҢ��}��o2�����ۜ�̈́��v��!�1���AF�� |3{���K��|�wbxx?��ϋ�.z�M7݄G}t��^N��9/4a�i��J
���p���#��?���������(�ńcn��&�K�j	�=��+�D��S����T�n:��00&�d���XNށ&_uY��{�l�J��:�b=.��t���/~�6m¾}��U"&-+2Dg�jM�CYc@ 6=���6�/�Î�1���NEc)�r!jq�}�9��T��	wv���c�Z�g��2��fހ�5˝���lڞ�(fL�p�5߬��v�ک^����:Oz3�b��ly*�j���_���w%s��Ї���T��ճ������W@�7/��&q,}p1��\��p)O�"9C!�ϝi��hRΧ�݆b��Fl���G�-1#CY�|�����z�,c-d
V �����癎�.�j�Р3y`؋�}12\�GD��eq�(������~FciX�ׯ�[�����e�{���k�����<tn,��Pl~+IK�-�?�	����!��q���s��;s�Ϯ�Ϧ�!#�j-o/��h������X�$�x2��ϫ�N �\5�+�\�AQUmNcsIPk�)T�m.>�d�r�5�Ϲ��SiFUm�R�lLE��?��p��x0E	K,T�vK�e��P{��J�-&]w;Bx�r�5�p��H.�31��W���fAǘ������Ύ6l�� 셃�Y�x~�^EDY��lP'|hK���D��%��� �~�X�J�V�K�����c�l�|�7��E��>�����˰�8���lW֬IC����𣧺�ozTy�%���j{i�wo��X ��¥d�tԲ-����=tN���{�2�����۰I9�1	�j�KE��	���`ݖ{V��:l7_��~���1�v�:�rYc��e7JJ�H9ȁ����X�ؾm���'o���3e�"�VX���2a\����l�d���g��h���bM��m+��W���_�]U�ƶ-X��^�D��J��,�2�@��k{E&ZJ���FV汶�ag��������s$�m�H���9����r��S�3����)��S�^��}#J�����'t��� e~v[w��t3�����v�~q��m,�a�u���*�&7����G��a�6v�s�A�dLJ�gfO$��5r�#�Q[�1|��Q�ǐ��H4���p.n��.L�hF�6��k9��_�A��q�V��z�uf�'}��l��,Cs�!Tׯ��U��J���*Fч��	����K�İ*q ��г��܉��v�	E�>]|gGF�R�]�����u�q3�DH�_V��?<�ӣ��5���%m��^բ�����Ѳ�6T�DT�Cj���w��ρ�`������n��n�C1ČH<�s3~�kQ'���k���~ǉF{QE<s��:�1:JC�!�L[���6<��/�C8J�Z�0ǁH9�6	��HH�1�I�K�nͨd��()�<�
�K�5�����w������qZ��}2|//Eױ�_���ɒ�j�'#�:�,k�tw�bk�׫~ȼ��Ϩ�#�4B����y�P���K�tȒ�T	�S�n���Z�����c0��x�+�� =ߴ�:/CX}�'=��f�6������Q$n{y�ReW��d%C�+ѧ	c\j����]u�#�Cs
�?0�̸p��/��I�������)�Stڱ^�ڔ���Ѵ��iTd�Dz�w�It�J��,
E=8����I����x��P{$v��!�tf�^�g7���+�<u]��Gz���Ԇ�T������\.IIO�<x7h��z���aei�<s�Z�m�4�j;��F�h>�*j��⫞6x���£g����p�Qb4����uU�����d��L�E�:e��+�V���5�4~���[[�v�G�#C���Qye�\
���q�#�]l��pU��(9U�l��[>�\�	ܗ��?��e&0��ZV��3�ɖ�g�]T��2b�>�#S�zl�z��9X����8<8����詯V4|&���Q�nQ��$���)e���f�Eo)	�	���`V�s�ҎQɶu��g��4e�K�J�s;zP[Q��>���s��>c,�}\'����-є��V�c]]�c]I��w�b+���)"9�����B[�Nly�bHs�ؚXN��h1�����z��3�\n3�a� h,�
�MH���lҷ]�}p��}\�Pu�H����^p_���~TZ�(US�^���ze.�mya/��Ӝ �b��&nB)�Xt��F��2��c���}tk7+�d;;f����K��*!3�+fX&3���L���oՕ��ѮV����DJh�G4�GM�\ e�3V�
P�t��d9v�U��F��e��Ҕ3kfY�>|�(&ٳ��$jc�����L@�j��j���Ud
u(q$�5�
��9�8�؈C��5���^6qX�6�#A��W�/L��?ލ���ׇ�C?F���PQY�A�&b�=���O�P�@g�&��u��A�`�c����^���Ub
�zϟ�"M��[&�1\|�4^�Ԡsb �������y�^\9�*�Nx��g����X��e~=�F8�*]��(Mb����uXj�f'�^���;���6M�:�άNrj3�W�}�S$c��{G��g�zE�8�%�S8w�I_#>�;���O��Z�!��8.3���Eh?/��Hʆ��l��H��k9�9��DʬĒfMh���ݝ��
|�f\�k�St e p�]�RH�P�B6�B����ԗ���x��uY�F��+�`�W�\$�Ơ/�~oH۳o���"3������c���r���n��}U6���T���Pq�u���63�1�)�YՀ$��r�/R��n����F���
b
��}����3E�w����=���=������Ug��f�>V�)z;�}�]�����	q�Ãz[F�;����AUU��`�WOS^��~1C��ߢ���˽�a��mӰcF����������W��']>tt�@]�1{��!��ߋ�	F%����2�D�Q4&,���}����9�~�Lѻ 8	�=��s��{{���p/ܵ�b1z�.c�w�����jf��\NkKb��Ӌ�7<������ΟT�v��qo|C)��"������	�	7�g-����1�f�C�2�"�0��F�6u���Wr��Q�}����U� v��%�����^"\WV�"����$.U޺cf[�n��Mݲ�[$F�P���I��]��.�O�]%����G�/���V�b-ҊbY4f�c�L�m��Ռ���H��ַc�소���5w*4�r*��c��]Uׁ�5۰�wR�Q���Z�pմ���� =��
���*�	�%&T(���dW�)z�_{�����}��)�'|2I��[G�[w�D(�h�EHj5P�:����*��jE���\ e�����f: �t����V�d��W�u�&��ʠ���k�kYJ���},�)��?:~Q�x�R��p�O�Q�J�^H�-
ӛ����Ci;<��о�X,VI�phP���D"_����Vua2���X';~)��3���P�<��K� Lgr��r^�o��
oڌ����o�)�Ks������3R�5H�ݨ�'�Q~�5to�55�i�-�}g0pi�lJ�D�ָC��mM�:ᙖ�I��1CK0��A|า:��GtZZ���Xچ��8ۀ��(uh{{��I\<���{�?�2H�\z�߀ϞQ�\u�h�����˾R�:5hu1��YlM	G�Ɋ�E�Kuf0ӧ?Ňi,��,"S0�H�J��U�d_ĉ:s
�S/"0q	�V�;a�wx|O������^~p0Z!%�7G�hzC+&�b�z�"u�,b�u��Ŋ���|����)�=��� WY}M=��}QN+1Nѭ���l�N���A�@��|T�DZ10�3B'��Ja<k���-�Jʋ-+;h4i9�w���ae�>���y4z��s�11���t�A���e�(����U�<������Y}y��Kv����`�C��FUV��"ӽ}E�}B��E�ď�fdS�w�s3�j攼�c���!leЙ���7�!��U�f)��a�^h=��lX҆Zx(&d�7���|(��3c�b��+�G� P=�ݸ���  n(�������;�[��MӢ�������Tb�r��ʔ����J���0J�9!���!�'c]Zc�=�ϻ��U[����ط"�Ğ��x���K�ja���#���mqUH�;�}ؘ�Bf��/�z��dZ�~��\�נ��S����=��z�׀����l��W3�m؉��?���Bo�:����2Y��Oy�̷��mkĢ f"+�2`�ޒ����)+eFn����D���{�Cx��Ö���kg��l�����x�e��x����h�ޣ�Tg}�0�"(Ґؒ�Ծ��8n��	e���oym�l�@~����bʏ>xLY!3���o�*@��xR@A�����	���s�b�.�b�"d-J��ݬ$� n
��3��۔Ψi��٦�s�hn`U۴���i&��O=��-u�R�I�Bk���W����R>@L)2�^Ō���3�K[�X���D�͊ku�j�z���[��^Bܖ��ʎ��.�RLE�eD�ԇ5ϓ��+�u�w�m�h/�_V1�����1�*���a�\H&���{�}�M�s���܃�z��J��^�@;7W�FÅ���
x���$3�
@ʝM��7��wL���P���D{g�
S��L�r��KW;�����n� �$�g�
j�Mu|a�2ū��-s��+l����'�ҾY��ӆ>߄ )��g5 e�o�Z�"�X[�����T�o��f至��̠� �:�J�d�Ʉ-W�UӅچvT:5h�|΀��s�?����⹊�����j��c?C$8! �&�YjPG.��#�a�nՊ��=}E�M�sc>�2�=�	�_Ly����s���E�|����qSG��rz�'�B�u��߇�c��ҹ2�>�\9��}v�N�ϭ����@�rT��5�����$�S/Ë�VD������.��o�=�]o�\f胢�m	��5ؼd5͌�����&�5�&*�F�N'���Q7�F\�#9�J�Ͱ��N٬�����������h�J��bJ^K\_f��Qס�F��Y4g���xY�n����Wy�y
g�N��^\  ���Xm����y혱����9�T,��~E@��;H�j1�:3c���� �l^�y�㑿>u��k͔9̸~(z}�NI��`) e������4�Ld삊Q
}��Ҷ�˯.Nֵb���2�̔�[u�x!��@�z͆,�Q��]�?����4�\u�[t(�Ao`�q.>��A�V�����c��^�r��KpS���|c� 3z�Q<\9�.W)\�	�x��8����&�xF�!�d�<��oh�Ɔ]�D��^�v��ϼ��3���Vi�b�Hn�F��C�־�Ɠ<�\'fX��y��fIK\�q|x�m�%��Al\�k�܋{��;����Qz�"��i+��Y,���̇�UVl��s��V�5��;>�t2�{��V��ɔPC'��!+��w�I�*x��u�������$�:���R��n Ʋ����a�[>���l�����'���R���F4�-���z�zz[4�c��u;en�Bْ��E���5h�]����1����+����7K���d�O�� �!S�
+e1�\g�a�}Qr�X��ڥT WHc�N-��� Rv���ܱ�_�[�*�ܬ�|�p�j9U����p��  ���[L��R9>4�-M��%����u��]�)י���\���A�I�@k�)��IH;�z:�k�^�0�(��A�E0�Pp�h�d��Q����2��M��>�c��pT�Ο��#� �|\7p̅��~XSm�_4!�V^���!�0!��#�@MC�\�(�#�5
�r��k�L�R�5&'v��T_�o�a�D"���p)nC Ch�,܎������H���1�ܯ���=5[��i+@ʷL)S����4m	�\ӸN�[S�Q���p�1�G�<(�@S�`̉��l�A��{�j*����/��P��l��|Ѹ��L��2|F;��^�)j�����-�]w?������!��kCO��|(Ë�Zt��`�����,?%���g_�O�b�s��Y����Y9���~�r����h �C<�Wr���j�ӓ�K��c ��x߰|ɔ�ĝ�ȗ;�;�"i�-�C�ۗ����4$�Pʆoy[�k��]8�"�B���mx6�,�7���$�e��e���≩�0�q�7�@,k@sIF�����D?��쉬p�o��7:#��a�ro��h�ڬZ�e)}1�n�BkmK�����<��^:�l`U�'�e0?@"����4�>�yL�D9�L�^�D�5�?Ĝ_Ӿ�_�1U���h/����A_�Zl�'g�Oۛ���lnVG3�]=�i5FV�$��U������w�h�9����^=|C�q�)+���ņ�-�,�d
��\ح��.�zx��\�T~v�Y�1@���Jv�R~�Ý{�񦲹U	����aS��ɀ�Ю���_�Y��ϸ��2Y����������4|B��.SJ�Ɍ���5o�PJ���
�8|������R<+��@�,��̠i�Ж5bY�y��Y���c
I#����o�gv�`\9��D��"h6��c�ϟ�'G<�_r���7H�ڲR<����?E�]e)��=�����¿��ݲ��~�Ox����n�G���l>K��cI���	�yT��Ns�W�csi.G�L�qe8�v�Hu�wCx�5�{�S��t�rd���!�:i?����uO�Xb���o���������.�޽Hp1���R�Yf�"K-f1_8{��_�=i8p�r�t�a�����A�L��g�T^r3���}�������g�c��~z�����=x����qebS�2y���t	���s;�_��Ƕ7�n}��&���;��c/�=4"!x]�C�Й۝1l��WP���e(B��^��JW^��MN���F9�;�<�k��.�8tfI�K����V����}xt�Z����⿾�_v��$�'���Aʵ��:��C��b��f�6�Lf�y�"�y�W��uRA��}�y�w�n� ��}�L.yø�9�͵e�q�a�W�5�7����W��A�WNE{9	����Բ5��;J*e!��	�۱�vl�>^g5�ey3LPj��1����YN4��M]�Pb�[����[wsG�݊\!,I��O���Z�+�O�{{�%w�
C��t4�5�O��m�2�o��"���:��^EO�N\���cS�;�3���XB뚏�TMl��+a(��:�5��މ���q<�!����-�p5ʇ����YlMX�,W��e?�@�(������K�{��7�yÄ�����E\ڄ('����ch@Z���b3��x!mWh�� �x<���ާ��-������T�g�WW�Gz�0����_Zp�P1�	J1L����58uɇr%��uT$]u�0V��a���ڒ'R�T*,�I�Y�=���˙�LƑfy��2)nnh����]yp��y��V��iI�۲%���q0`;�i!G���t�L��@�N;�%%L�@��@���f:@&!)�6q�����6�2�й��]+�n����Z����dO�̼��c�����}��}^�H�t��}�,Pm$o~E��%�����*���7�:��^������"H}�]�{��Ú-�<�3�㟞8�}�5���3"��x}��.���n!ru�-��?�S��M�zev�M/�a��k�%j�]8ٺї����Z�i��NV*���Bw�����,�~�v�,�O�[�C����rh�a�������B�V���(�-�<f�&���/�w1BbS[U���a%n}g�(@��e���4ʗ�ӠE ���\��|���B���^v�6"���Q�����+�}>\�{M'ph��~��+�\*��y���[�������b�EJ1�:����,�,ǉ+�
���^β3�Ch��&��ơʾ��*@�r�#r��>8�k�Z�99y�ۑ�a4|�&���B��3C�N�b�9�bܭ8Ϡ[4�j�:�v��݆���p�_�5ř�rn*����ht��f�+6W�bIp]�>�,������g�:<&06A� �ٽ�v�#J�����ӱ���wM�8�Q�U"��xZ��y7�=�l��5܅~{&��\�\�W���#8�Q���B5zcg�ZW�s�z�_��{:���:ԋ6�����;��{���7���w �r�+X��/�`�E�PN0�߆Q�Y��WcLQ�^��Jۧ�Vb�� Vt�W#�s"'G��8�����]����F�����VWh}��m���aDb$#H h\$���AW���i�Є=jq���)�z9zO&k}F��L��v��|ۤ�Π�#�$8ۤ��	vr3�6�)8+g���L�Sv�o�r�U�2��͡B\�R��u�[��}981�R�턅�iο1\,+oeD�"�D��j"<��ن�r�<9.Z�U�HR󍩬�T�9�G8q4��f�>4�S$��b�G�wR���:�o�9��n���q�L4�����H搴�F���H��#GT7�}V �@���k�d
�����Ao�\zT��TK��u�E������T���M��x�����M�[�'UO���Z)��#�S���s~�(�4�>�ͮ�l\6��.�i8�ܨF�9&��=��Ry!5Ւ�Z�=%=^� �)����י�"\���o���<:Yg�>�s���W{���*�2��8�Ӫ2�h?���oFIf���Z��}���`��E��qP5���A,Ms@�a��{0*�(O����E_?nط;�l���-�e��&����kIi�=���"�o�B�G���xщCf�r@���R�0��FM����AeƘ�8��;>����p��k�sE.�D'#
;�{/�\�I�f�%�ıX`wd਌�sԡ&d?�Q(Hs�\��ъlȹ2�jeВ6~��=K�C�}�Eؾs'��b+���L�R���̬l�9�Q,�� ��L�/*4��
��.�2kw� vd��(ï���q�x���x�ָ*w �����kP�|c��F3�\<�U�#�i��\�1nپ6윫))��E�Ox�v���!-��x�	��L�b�֭ؾ}���s ����&��1�q��������yΌ�ЫLی��P5��B7��F��f�ʬ!��Ƕ��nkYی���Q|��[�]����Z�Ҫ�B�M�~�>1�����|����-M������S�`�`�ħ��f�o�EŒ���]�|2z����>��]}ʖֆ���t5o���՚}Y�Kk|����k�j1�G�N0�WqVo��_�1o!|"4��Ng
Y�I�/�.����l$�b4��EK�'�#��k�u�:s��.mt.�Z[S�]�b�,�^Zc�cT��n�YZ�k�]��D��u��/�J]��)��ʠL]'�6'g���f�/-<#��k�n�P��-h��ҌI�2����1� 7�5���ԍ�Y��yvfi5C	 3�6��KFF7��[V�d�²g��Tx��E �eɣa��'1���/n��ӷ݈o���ۚ�:e�-�sm�ǓV�5���Bog�R&�2���NR��v7�w̯ˤ�b���sZ�@�9��U�A�� �%!�3�m���|��'�H�Bn�DB�Dӻ��5P�(3����6��5�*���׭�ҍ��p��24v��V/2c��Ԭ* ^�w�\�ϾHo/z��5:��_wT��n��WX���v�7���Q��z{�ƾg���1��=q�=��Cݓ�B��r��p%� CCC8r��H_h���뮻�m䄑d �� ��7(#���L��*���m�H�� 5B�$�
^��O�ѵ�WlVe����4�?�����IT���������w�Wym����'�۞4+AYn����~]���z����Z���mx������ۃ�JY!{r��46����e��|�ǲ����-����5!#X�k6W���{��U{Y�������D��!x�%t]D~Q��Ɓ���������ٱ��oʏ;'3p���M��K�;aӍs�����ܰ�
?<|R�X�0˩��(��%PQi4Ӊ�0QD�����0�XH0�y�����ڼFӔ ���s(�3j�KOl<׻����[W�Ye�n������fx{y���\݄�SqDL|_��o��sǽ�n�6��Ki�R����*锠�	뤪��>�X� ��6�+��fK�E 9.�z���;�ke�it[�_`��.Բ��i~=��HlRo���r��ru����=��[�7�0�m��|h8�`��H ������2��<I��^�����XV&�J �/�z�E��[�S؍g$a
3)a���H���'�/�s5��ʤ�� ^��!a�]���"��V��
T� �#�z���% ��Du��F�d�&qQW6�K�{�E�₨y:[��3�����B0�z�!�P��� �^FPÞq�k�c[�Pf�
)7�rpz�`Fɒi��j�n-lEma��V��æ�-]㥁2�X���R�}�zT��i���n8E5d�U���3����`6]c����|Q��������VC��G������.���d�>���gݍx��MbrLS{��}RKkl_�v܄�lk�h@L��~���j!3�"���t�_W����;���z����m��ΡT�N�[�@}bX����K�l��:�^��vj�O����!8N��tUn*�C�w`wv֔`��k�������r�U���3ޓ��h�Kg.���R����7C�k�a
It��縃A�	)�Iy�TS�d"Y3��ŀٟۅ+6�f�^���
!B�:��|=������W�{�9aK}�se�v�����`����%�NTTo���C�}=��A�DL����74-�0��Αe����֖�x�=SVV6g�6���������؍�(��`�s�U����>�A���YT,�6��_M�,MG��cˑ.1Y\�l�Ṕ[��O���ە =�Q��z��&պX�YB�ܱc����̍R����?����9�R��"��7��kBc�I�P��|��Չ̴����)�A-�^܁�63�W�HY�7�v2շheR&03�������q�2;�/�\��9s=�DH%�����i$>�cP 3eܖ�p;�V�V�L�-���nF�d�&�O���Jw=�ZΣ��YY��0��wF�����Hvh]\@�Y�s�F�.����R�Ő!LP�%qg��9m�����aY\7��e���E���安"�!ZVk��85Z���2���� ���E��d:���A�#8�хׇ��!хr�z�?�/�r���J�BP�D���k�T��L�����.J���qR���P	V:��v�'��݃��%mm�������[2��)�}�'{���:�d�م�fp���/��]��ﵩ������d�7j\�L� _�J
����Qcb��3�lj���9�<&ˊ�l��T�l2@A����̜��4Y�6`������I�YK�]Q���Ƣ<�ٿ�T��N��_�J��4���������a� t���/Kq�[�2.���;Y��#<���{�~�ӛ0>a�y��Td;�� +\DxAD�Ud���M�R0����ĉ*�w�ܩ�&2��=�v�
�6��� VMM���oM�y� >�����ǯ����:|���زe**� �566��߰aCX{��*ǁ}�9q�]�c���*��[dG$>~*�C��N8��e�S.�&�;�f�G򔘅�i��O:�ʋO�G����ÿ�g�j��OW���E��*�(
%�Ya���>��F�~�i��W��v���Q��3Ϡ��ZG/�O$S�]�jՌ٣�a�����E�����+���{�w�y�>����s����#�<&��3+K�9�
a�3ٰ�<|���^�||8�5�}?`Ǆ��,�>R/��5<������9b���3!(3ΰ�HDr�e��8Z��y��D��bB`Xg����oy-���<�\���^��Au���Α���$\�4����	`#�KKK��k��"	����=/��,�/.AX�Y]eX ��&��`TY�611!p�� $�\�9>9�;�Qc)�uC,D�F�w���E�ji_���ٳ��`�'#�˄	ΐO��g�<#�Ҙ�E�o����E�M��J�S`�8#�/�} �I\"0�^*�====J�� Fsf���ҫ�B���_2'#	B�ub�f&�Է<%�Fi7�G�2��U�q�'�v�?���%��A[HY��#J\��4f�S4L#�+�:ǐ�L�0������o�|�D�قU�`\g		���$��\	b�?��Y���c��O���Q>V�vg7e
q'�G�c��Ĉ��k��i���\\� Dp*�=409�LZ�%�f�7����ރ��@o4DD���y�������+i᧕�G�q�'�C�K΢&Z��O��!̖���AZ�-����px}�}#�]�h�z9�YI'��MZ*��\��1�O�����>ĭ�aB�FsI�U���7<����yi���j!M���u*��E6w���ۤ� �E�Q�e�|�9�V{�!����4Ї"��%p�����1���)0�4�=%��+H�Hgc<0�ԜU���(���Xn�q��v��r�$@�='���H~�+�lND"�'��#o�e~E�-���{�X���؈(q-cL�]��^��Ƅ|��n�M�6�3��X(��+���3����E?��W[[���v�]�vzDOڐШe<�Dc}���oN�(��c��N0� �`�s-,v5�Dx�v���<�܍�[Y�!�hd���y�*q�1G�ƍ��SO���qMΐhGd,0���&Hy?�����~;n������}��:��t�k�g�)-C��M��
��$+fG|~W�s�?�2�"](��D�K��"�"'A��TҀ�}�QC��^Þ={�nݺ0q�	�o)�r~$}��n���ٌ����a����@��ov>�i��'&�ym�jݸΖW_}5&["AȊ�ĸ�٢�]]]��r���+�����L�;v�y6+=��|����('7mX�����Hnmm����!rA�DC5�j,^knn��Ç5J/�n��__�L�M���xg@��|����/��X����=p� �x�pNs/y5��"�Sq��]���E ;�]�w�x��򗿜�pT#4=���g��-W��x����g?�H��U�b�_ ��y~~~~R�׬ĺ�k4Vnf �tP�Z�f��p�'J7����� ��rd߾}ػw�a$�wܡ�Rq����~���l�-�ܢ-:�$\���j�����&OG���O����p�f�\"���/3�J�Kau�e ����$�]�,�^���*�,2H��o]��.���)�xH�X>��]�f�*E�P16�X���C޿"    IEND�B`�PK   �zxX;��d  �)  /   images/35440911-0bff-4ebf-83cc-bd2192eee111.png�iT�׺�7�RE��d�Q��J@��֣�S�� `S�`k� ��=(�ZE$"C$�2�HB�L	$� !2$���#�ow�u?�{N�]��o���g����#^�W�X� ���w���`	�e�"�ƕ�?K�w{��,KGqr)��<�;? �<Q�j|��/ ����},1o�W�K��Q�dܨ�<��銗�z�~�ƣ���޳��kwuo.9���-Ƥ�W�~{m�}�}�'�ﮤ{�hK����|É��ܬ��
׵�&�1L�^��>sN9;<�/�c ���6<7\�����;�s�t@�g�*��	
f�l ���������2-�ٗ* ~�d�d�d�d�d�d�d�d�d���&��v�m:t�nQ֔�St��&�\�}>[�[W�����<���ek�]��I�\���3�ax��Q��;�>�sc�gr�Y���=I��$�1z�!K�}I���z3�>L+���	�څyʂ? �}�U?�����v��&�Ρ7PCϯ��^nO�p�<�D�}N�g��Q�(��T�"��%K[��9>�yUot�~�Xs�"��z��nX��P�G��&w���{���b�4u�� �����	DTOs�Я{��؁���cn�3�|��]~.��ϖ�������އ�1���U�n��U�Aoѣ[R��f~~~x�A��y��ۧ�.��v�<e�&"eۇ/q�o��l�o�	�}��l�4t]���0�B���9f��]/~A�$hE����L�5e m%_��4�E�v5GL�U�Q�C���5�:NTZE��H�o�~$���<xyN�CRiNyzhSF�A�ꊉǂk������p.�S�Ip�쉞�~W)"��5c^��q)��!�Y�M�s��G���(�Ƨږ.�it6<N��m�6k�g�����E��{��}jԗQ�t_P&h��Z	ƿT��r���;`E8�b_���Bb�|����R������9c��A�ۗ,�#P]%����#�-���H�ƠM��K����t��JQ�T)X��D��+�h��\��V4�f���1E��pf�%��n3E�� �|��b'��ǯF��[2p/;�����N8Rל�XQ�Rj�0�U���#�1O4�(��S��>%}'�;�mk
�M�Ǳ�A�БQ�;ۋf0��i	��P��s� �i�Mhz����o�<�q?����]�+�3�R��7ۦ�1�r�AA�G#�� i_��8�S�`&�y�|)���>4��N��,��ܤ�2aܩ�����ƶЦNKe�嚀��j���D&#P]�A�2��f�����A{�('�KG�D�p#��K�8/M@�O�i�閒l�_� n�&�x(j���ޜ)4w��Q�y��j_���my!1��1I�N�m?�ҥ ���̓4[���O3U��ʉ����	L������v�C�G�b;P�\��tX�*q���&`���{�'H�����ZCIܻ-��!<hk�7ǋ�;�ߞ���]�v��s�{� #n���i?u��
9�H�s�bC�O�7�k[�(���2�c@��+;"J���6]��>�]T�g��=�VO����d�:B������u�q��������,�Y\S����=�E'"P��^��FՔ��-��"@\�Oq�$� ��� M���r��B�s�W[(Im[�Q��k|� �,�H��?���=�F�l2�F��+�q�����mW�]�g��f;�ý�Nj��v��ɳdY!���BU��:w
�܃�.��0�:k�E���Im���d�mQ]��й/e"1��${��Ēf��+�q`WBD��Կ������>���'�Q;q-������A0x�p%˳���GC=\���NO�����i��T��:���m��}'Z���=���w�`k�+�$�'krt�������SS]��F�K��_�T��TE&��(���c -d�e���Z�u���P�ry��{�Ly'������`� �K�̼�dQi��X���@k�����;��ӟJ�b<ð�'�@4�����U���4#I��r8�d�γ?n{L���SB$�(&���K�\g:C&Sf�Q����v5#C%��ر��.���&��mks�I5�P#�y��'��E`pS���2�۾ט#�-��/,{��,��E
E�[)C�9+d�־�ahh@
rP�"�:ɯ���c5��z���4
�=y4��I#��蒨*IWV6�V�ۖl8��>�쇧X�m��hwZ⻉�)&��&�M��#{���E��B��8O<��6��}���|)��&�����w��؟�^�4��Äm�8UJ_
���c�F=^�>��!��7V�̳����զ�̽�Fl[����O��le�.g0T"�q	{����-v�%�
�>.t��w/��΂j#���#h�_�V&c�ͳ)���B�M�e
9c��7$>�0T�J��|5��f��PKg��r0�&�bZ�]5IS�b�-�Z}ܱ?�;(�ݽgz��C�Z���KH��a�z���F4\6�#B�X�_��ۂ]���d�^/�BS�DK�3o�e�����7{��A;e��B�`�2#|^�8j����^�1@�O�z�*9�_�B#�E�jFk�4e�?p��	��q�^/v�,X\qؗ��!�HXi*{F���S	�_����fdOE�e�m�
�.�+��m�����M�AQ�3����m��{vg/��o�4��$�����O�P�n��	�Ҵ���ɓO�E�<���Â��'��'�_�@2�w��cl[�J��D�� ��!�]�R�C�a��`�!R�+r��=a[�-�Hd��$�F�|�j~=��=d�S2��nK{|����l��ո��t�M͋(����t%�_���0��yK#�}����Q'2�o�AuB��?�u������̎���K	�c��'Z��	*/5`ZJ��Et?z[ynή�0~�CȰ�}ܖ�䚳S��LS_JR�"Uqz��a�þ,o(�T��bQ�S�il������A�B�y�����?5:H��/#��r���h����B�d�d��eB_�\�(��w�pӡ)�݅�=��qH-���7�n�3UwH(���M�R�{J�k�}J�]'���gf>���a2��u&�
�����v#�īO
U���iw��U�����	�hB$:������k���Zon�k��9,7�������S��M���~�A}�����h�3��:(�Q�W���f��zuY��,�#�����Ab������K��I�A���b���	5p-sǻ?oD��I(;�V��FU�(����8l!s�Ѻ�q����b���:R��Y���؍����P�_��߅��G(�QJ�_�A]1ڹۊ�tUr��55�g�pלF�{M�c^mc��de��ᆹ ���Q������W��gI����f��|�[#����{L7�a'���S�q�w��Ϗ�z[�'�T�Ǻ˝�M��aj8m'���:�=��o &��SrR�S-��Pt���k�t�iK��:g{Jk4S�.$��SRgH��)>�x��~HM���PuY@P��eG¦��W�n��\���n��x�u1'�%V�].]�U��=�ICG�<��Ԑ�$��\�Q�]'�Q�|�>�c���A���������1ϖù4��H�D�q���mX���nv�>$G�8�9��(l�S���ǫ�T��}I�@[n�@\����X���{�t+�uZy�p)W2jEa�z��mp~�;Xw.i*�ܕ"G�f�]|�_0CN Y�ʵ�Ou�6��ָ���'��u*悵�A�߶�r}^� ʫx�r�[��}/O��	n������������PՅ{�\�5p#{)��^��!-���'t�}������x���-U%B�sKŀ�h�v�c�΍��	:ړ�Vkb��Ǎ���O�;�͗����>0��Z��Vd.�i)J��M�s���[ơ� =*��J���5j�n�o|ה�6h%Y8���ule���-E"�E��u�>�2XJ�`�rk�����El�c��ADH��{�zf|�����{DR���_��;���葩�`�)���ǡd"$-�p�|��@h<��
0ރ~��V�%�+2j�i4N>��Q�����D��5���ua�'�0�	j��Y��<<C�+lK3Asw���nK��#�:g2����U�}����N\�pH�R�|u=��R����4�t�#�+)�5�5�+Dhxp�������uPNlP�����,rG����BTY�����]��+)���4vCTse�d2��c�E�?�R�����H�j/A
�'�k�}�?�ۦA�Ь���0}x�/oo�<W �=�Q��Ջ��R��p�����f�o�s�WmwQ�r4���e��gD��Ǳ�m��cC�,�qʾsS63��W�����F��_D������{wV��p}�s*��,
9mPU�Ȏe|9��"e��g�a$d�m���6���E�񊎫��cyNbmTHg(<��U���}����l�G}e�a�4t�q@Ε�Y��j��u|4�~�W͙)� Lk�LY�8T���X�=sG�Id�=�J7ռ\.�jM~�l��3���@��d]��h�7��ބ�w^Xnx�]qa�2@Cz(�0)G^��G&}���i�f�҂��Tk��e@
6�;E�@�Y]�dԹ-̱8��Ġȝ�����G��)d���&�z�:�(yo�������W��?��Y$ϞT�xzv����h�f���m�+?�&�v���0$� >�Ҟ�����N�W�)IQ�Bwe�"0ҥ�J��ј��{m�s1�g�V1m�N:
��Tٗ*7' q�T�B&i��]�����~�J��3'��i�R�m�����uQ�z�є]f��F,r�w��"m0]%��쏖O1��yW�`��
$�j���^Z��F}����Cj����|)d˕:uq5(�^aEb1���k��I�VS[z+ˣf跃0K*.�p�a<y���l�g-���~�K��&�*9lPz��Y�L�ϧ3d-�Z�T��j�b����~Jv�31����5�������p'�s���c@�Cv/g��clڼ��
%oA�J Ý�Du�<���~^�0��k���-�*"e��:��q77z����wo'�Z �7��ӄs���I���{�PQ��B��0���㕜��S)��݊��ҍR��������'���+>�\}
3]D�if�*#� uC$-�1������kf~��O#������b8�7�e!�~�`1�!S��Ddһ�Bvř�~�vf�N}S��܋fԂ�@�8̿,dox`\{#���J&�x������ �r�>�;�Uկuuu��G-Nww꼹0���uhX3��ũl�N��ۗP�m�8~�3g�;ܞ�ֺc�I+�H���v�z8߿*2i����L�j�J?�e���c�%�"��d��I�q�
-C�*2���>�Vʃ�<��C���Σ���Zk���v1�2��'����Gٶ8�-[;a�ۥ/��
�� ��O�����E�??l�4�������<5�.'*K�[}��%�֮�*���p;f�!g��.��d��?�mΙ1�	��5�2=\�w'��}�R."D6]$iEJ�q�;��6ubL�ظ?tYp����W��&؀���
���9��m	G�9��˃��?�PK   $xX����+  J  /   images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.png�WW0 �]-�+D��DM6DKV�Ѣ����Al"�Z���$z����:��V!z�������g�=3w���=�:Z*T��  ����[��E6ٝ�L]�{K@OUco ��� �����|�`>z>k/{ ����x�Z{�xx9��J=  @Sj�r�o3v́�I�L��S�g@`
�\���EG�T<e!�����DʲϘ��|���E-	:3עt�&^7Cx�-��
H%TH��!�U����������C��ח��(���~�|����>��`����e�~�L����E`"#�n�����bng��0�d�w��f��u���R?	X_�B����������`؂v�r��I���ӑ1��ԙ��*3~��_��:a���skZ8��[;��"���� ���p�HZ�������1�d���g/ǚxx���L�	K��%y&�Zt�Q�� PKI�!����O�Z��k�>)�|yX@8ҳ�́ߖ�N��+a�i��?���m�ޢ�[e�O�M�����"si�n�4{f�g��!l�4eqz� 4W �J��(����3=�ͤ�;[AI=�� �Z�G�'�Ci�55���T�eqo�Z�K��T���/���m�p��&�5��(��sց�ѽ��;�:���v��F3��� 氉2��G�;H��1��"�{I6WY�#�JJJZZo����gKJ]����p�Y�*�`��&���i��&�k}pp���F�oʡ�t ���>�x���n�3c�ºk�����Vq�[˛���ai�ɢ�L�7~@�ĩb5�W����`S�O�=�\"�����j��oq[��Z�ޛ��~z�G��/��G��)����Ci�h�k����i{(z��_�zģҕSD�i�����SO���"҉5\�^QY�u��6W-"RoMaJ�`:��󸼝�@�&�GH(��3wkװH<2�wgv�9���>�M(�Ѱܢ�k	u��WKJN>��`�i�꒬����Bfxn'�R��c`P1o�9��T��E̵��h�ޑ�OZO��F~��nL,"�h��UO�����`�}�p�P$v�"%Ʈ�Y7;�>��B��Q�2��'�З��>Q���ߨ�|��>SU &N	�}�C��<&�uDi�ƴ'�5_��i��H��dƱ\�7�[�i�^�6WŊ6G�M*U����o�c|��3��g��4jf4�퀋�Da���B�h�bs�H��Lu���_b}���p��9�ib�h�Hm���I���� ��w~�:�Ǚ��(�Z���iaa��-%�X�0n���4�S�P+ҙ=ߊ����D��BmvI�Mm>���}K��A�U���q���LyKHk&��MjB��}���A�f�)���D}�ü����{����h���xܞJ�tW�&P=�a�kw�m_,#����rׇ�߶<J��V�vg���^���ҵO4 ����l�IGB��L��PS��ڽ�����	�;m�y�}a�.��%\o�jͧ�g�# lF�<���s\RCj�ch.�5O</[ߖR�̔��{o�Zwu��H�UV�E���_�#>��N����1�+��Ġ�E٫�ͺ���vub��Vt���9c�M�j]�򏻏aj�(p$v&�99�r�ئ(��J��Y&躙l��u-�1�}x9��x�=Y��絗�<D���T͢Mxf6���Ȉo�����{�W�������fF��Oʁ�����w�7���C�f�<�{a��ḡ|̴n����*��V̶Q�$��e���YWc8���dO΍��$V� =�z�z��!�Nj��8�H|������~@�����;/4��ʽ}�Btnb��D��WsV�_዁�tPY"ۃ�t�����P��~/�9žcT��bQ�F���n�}kM�F=��(&�����<�{�W���i�1Ӣ3F\QJ�"�i3���%��1�ixjF��aƓ��r�*:H�s�Q�"�@�g�����������$-x��d�۴�D,hO$LDRS{�T����ib�7�G6CK/X���7�ɣ� �)��֚��tWDE��+�9��R�dV\�Ѽ����E���X�;+�[���P�a�Ze�J-s3�~v#sA�;~�sDh	.l�//��ܦ�:�S���Ż��|������ᬹ��FO�����h1 W�f�V��e%����\+C�p��T�8�wʄ1���l�5k�a6�|z��j��������2�zX��:�ϳ9	���P�������@�UlA��0Ԥ����\[j�4�r4�j:UOz����'y)c5�����;�u.S�����t�i��p�*y�0ؾT;bg2015A?�Wj�l��ۢ�$1ye��K�����E�^-����T0���8��� ��p��a
�`h*�Nj`���S�^N���dB�@#�*N�CK����9���R���૕V��v@cy�;�K��z/:�,Xi6S|��궣���M��v]�� &)��\�4���9h����_T����,��u��=�n2�O�R$گ�[?&̽�W���'����>�޸��R��q�ݐsW�t�)���9RqP�`��]�
� }5
B����g	k��g��wf�Hf�1bt��}����8��c�N,���.��)��֩LS ���5���梓EjP�r
|-�������q����F�(���5,�y@� g���Z WMP�;�,8#�]$.%'g�^��!��.�x-z�\��������NQ�{�zAz���Qr�����-wT�1�,T��r��5:}�R��`Ha�ځ_��K��������`��s7}��3���ڑ_�129kzV�0��� ;�#+w7�p�i���L������ xT{�^W(qm���_N@xGY׿�<�F�^�FNz079[WE�D����i5��n����a�Į<�={�ܕ���V�i���ܬ�K��$�GȰ��ץ8IU5�D:9��W�Ռ�,!���%l{)�8Do�P�H�~5(�\@��S�mmu�e�m�ڥs��>+��ڃ	:=s�Cl���Q�X�f	Ǒ�V��a�<Z�5#u&r8▴ ���c����~��?�j����Q�EB���C��C:��h��a��L�І������l�z,.���'1yiV���F?��K��.ϱ����"�lC�&A�{>�v݂���`Ԏ��:���<��Pj(_�q�e�E}��*Sy�ţ��)�E��k�����N>�a��Ȼ�U�Mċys|���_�֕�d�.#pѫ��4d1�&@�h�[�Q�����仚b.��W����M��R�k9�FY=�t�fn<O%����\j�l���t�r+�����Ñ��T�(E�@D�����3jbT��hy��b��A�`j	�\)�v0�	Ăl�r]�_��_�%K��*����d�PS���ſɅ�.��{ӕ�#�X���b�\6��K�g��,id�dQ7�o�|#�p���JN��w��
F�$L���2-x�s��`�
�,"#���ށ��1'Э��x>���
#����-�|a�M��^Zօ�Q����q��>��Ւ����v�Ur ,��[���t���(dN��z*�Vvq��}zR���j�fC�;<he>��4�d�R��f�Jso���|���_����|	.���۷�R1?����#�<=���	�of�d���{�-����k}2`Q�5�����/���q���w���t�B��a�˳� N��%y�{�es!}̰B�crY�	5C���ņ-5+z �!�K��U��9i��hE��������$M:a��Y�UmW���JU������R���)�\�Z�~[O��-#���b���T��\p�������O���h�_�fR��L�����WNs��B����z���{Xc"]���oMe�X-��sī�M�`��E������[���Y�T��0�:������ϟ?�=�
^p�>f��ݚ�4v1>�^���f��"ȴ0��^�f���J�j�M�ZŐS_B�M�/�������c;��[�sCT��#�܆���b���?PK   ��WǆO2K 9X /   images/59f150f1-5697-4080-b5dc-b8b306a70e65.png\{T�m-  ��)ݠ���(Jww��)1t��� ��twH7�Hw3p�������w�`X0�<�����{ވwo�1(0��j�t�6�P���4{�����*ƨv���Ro���0LQ���.
��/B�O�8����BE�����A��,����'^����E�=f�Ք�}��Jx$�&�����_��{����	����:�:��z��	�=�e.Xz���Ո^��HT���d��X�e4?qӜB��6���Ĳ܍uN��i<W̱s)���n+JJ��|�����H>���W��7.���,cr�����!������jS?m����߂�yW\ɇ���oq�+-���Aϗa�k�?�����wh����E���W<��R��\�� �-�}����o�o(s7j!��n�9��;��y�km~I��o*F�]��������
^_-9�\������t�{���H�Sg0JEQ�U�t�X*�oY{������w��ݶwO�j��9H�`�Gۑ~�����0\ڜ�۝\�J�vt�tƦ���Y���s�,���87�Ȟ���8ԯ�$���b����^���9��xas����	�A�)O&��H��s\OU�S0�i
��v�~��[�rԲ�����~��}�S���ʇ�f��澅���-?�+���o��]�S����!��7]Q�JWΊ����M̍���'����/�Aq�c���@�'b���bh%W�d��1¹�j����l�˵!mS���+���bZC�J�]�����v5����H�����/��J�f?	�gl�72.a���}S�ʢ��K�C�	_�=��g�aS����] ���ۘ���=��8�������>��x(��`ə�`�;� ���ظ2�$~|յ��[(Apy�
L�	-#�BM��&}c�6�t�����e-ݝ�>�r�mg����`���v��:ǧHt+�y�����B��[���{�ǐ#Eo'�(�d�>�YFg�Z��|��Zv�o6���v�E��\w����Q��!���l���u��p�iݨ��(���w����UԜ�E��791���V4~B��9a�~��sn�]Q?�͵�_L�{��{ָ{/S��^���25[�z��B��H��#֜�^�����i�8l�b�7���<��������d]�gl;�*ϻ~-�b�TN}�z��|��ӭ~m?�5�+J��jcӈ5�%��/O�r3oYM3�˰dL�z���Q�٦G�����v�8���nQ����'�`�η��u�4COW �O��F���%�d�Y^{\�#��@�3��Lݣ��8�*���g��d�p���vI�����l�席e�}\���#P�َ��+�6}��T�-A�C=�)�l�v��%@h��Z��<���aӚ�mwv3'ݥ*���|�������۳�����\����R}������	���h����P���a��_ss����̪9���i!U� qU�F�Q��]�x��|���tF^�4jya�)�jV�7IU����=�RV�`���)�Q#	~�W�K�?�?�1W$�,|a������r���re��-X$�Y��U��ͅ��<<�Hz���r8�Mʡ߈��T���������f�=I=\5�è�s�wP�|'aq�I�Y��/��kG��CH����÷ 
�lE�b"�e�E'��W�A�dF��ewŗ�@�V����~�Z���`|�T<N[+^-�j~�!	[� �E�'@��&���	5i�X�Ea�Z�:�����{���k��d4|�v޳<�oތ~Y��ƥvZ���G��Q���A���F??r��f�U���s�H��?����r�kA�2�K�|���ءs���q{ ����}b6(J�*�7#��a�˱���ȫ��TDC�D"�.��h��I83�Ŋ&�G L�ͥ6w��j;U���g�Z6�@�"����U�̩�p��6S��BjS
���@~2�t�����2Җ�1�R���T|������I�M�u��V��3�������n�0_,�J�j+꫟*C�[�
~\0.C��@���h��"ƪ8fdϩ��kƭާ��@9Z��Z�2��%���zUԎ�P*VE�s�gY���@Ŧ��W�'~ E!5q�sh��t���T�o�D��N��@oĤ��ԟv<���������}��DN�	�=owX(}�-`sAϲ#�zH���l�b�10��l��e��y�F����q�m�����`���� ���y��2 �q��c�Y�"�1���9⮛=�����I�~�3�U��-3﹮�(��Ҍ>{�a�A����ˁwՊ�(Ũ�׃,��5��F%ާ�ӿ9S�Z�D>#37ľE���Z7`�N�����Cz��D���%�a�Z�z���ruY���C�T���<B����!�7��ѣp�) 5�o�p���
ءEmim����O���(a8M]ə�;�E�������t�������a�@��M��#鼧 id���W�ъ���*�Q?�V+<�`�6.��i8ujr�2�����YZ;�}�lc̔��/���t�
� :��ϑu�P
i��)X�K! �����Tf�lϱ��Y(�L(��ȹ�p�W�Ⱦ(�����G��Y*.��#�-2x<�#��ǲ�<v�R�l�-ҝ�-�競1ԝ�Ls��gs���
��'��2�;X̓y6.�}���< YEI��b,�����`g�ݡ��ߝ��i��i?m�iww��Au�55>�R-�_/��D�e�k�将�^�I�u=��~c�,�N�EW��Ikg�[�=�����`\�2�����oY�5j)$5y��y��J�>���� l� ���q4�Z�(ؠ�oa6��q�1��!����kr�!|Ԩ�9�ںa	��*���4-_�̴������r�T��+�������K�Z%�)T&�x�T���f��e6��w�N�-������Fa�&�v
��������C�C���h�ޠ7�K�S���-(GА��`3煤���Z89�ڣ`%�	�۠�(����e��9
mr!#^���?�
8������"�N2*��z�48�okVٵ�� �R��;���K#5�_��tl���F%*K
>P[�$]c�ș������)���;��6����I�����v���8 :��� /��E�w���`�;A3����º��IV#��T�7�X��i�WVJv�e�[�x���|�|5)O�t�cfĒ���\i��3�uLd9��ދ{�W�1�؂�4���\��;-6��g̅>#�̥�a�[� uE����4�&��~�L�A����僨��Kw@l�U�4<ZE�5_�ڄ}W���y��$��?*϶vѺ�����p�F\z��N��'���rM�`�<2)����U��P%�Ի����-�WJ�<Fx��ܺnL��H\���ȓ���V�2S:�7�&��D%u��o3��@���Ń�~�F=�Q@9�&Lα�č慎ߙ�Ͻ^�M9����b)DRp6�R`5�~�@"��������Gk2o�9z�0�O�~�m^�����>��r,6[�3��C���#�c>���',�ʢ�5¬�h@�a%j����95��o�6x�d�l #���V��+v&7JP>~o��I�#�e���*G�2�������_o%�Q�~I,���V�JB&�]6�P�H88-7; �S�όcG��Q��������j
Ţ�mg�$��۱8��)�Ɏ D�����!�>T��~�����z9��rLk7W�-�x��BN�y�`�k1����7�
1er%F�7�h��F��UHbG��w��|��hw�T1�-ʒ�X�'�?p���r1%��]!�Ϙ���x�*���r7�d|����fPq�U�D�x����������tlW�����"����U%~�y�Se�4��)ؠ�%��%����B
�f��~A|�xA1PǎY�	��3i!g�r���xR�뽙(^MI���V_Li�Kw����E&�T}^����������ȼ�TW���n�Vhb������Z��
e9��vt�?Ò���^��q*���7+������Y#.h������8\�aEz��&	�T9���]����T���鑪L��4dz�1������-]*�s�f�����݊��I&�K8d�e<5>F�o�zj/**��G��"��jk�ƥ�V�^uDf��/?Kg�S�q	=,u0Ӓ��VV��Y��j<G����T���������Rjd�wU�[�y�p&� ���*b��U1�QO�:6�|~�L7!����F����5����D��dZVy�Cb�>5�ta� ��~�4x�� k�`~>}{����P������ǫ�S�e_N��Ms��Z���vO�ћ;a薓+�wzzy���Z�"���8tϾU�������KJ�@���wr�g5�Er���c_2�TsKc���<b;*!J��6��O�*�7��1t�{_��-$���~���x�%�K^�jk>�/�x�������yUz\Fvݎp�DK6���/Rc����X���{ޫO�%|!P��ѳ;&�2:�2���Pn�������N���;�P�°�Y47�m�Šʫ��2UEB{E��΋?DmJI�P(��S���	������)�=yZ�:��NĶЩ��Ɇ�_{���� 3y�;��V������j��H׀ܠ;.���(追�z��ݝ �5�q������}���ޞ��θ����_L@��	y�}w�C��(�d�1)�xK�y���'ꨶ�!u�&c �j���'�~<�|�r���w��2`��Pq�^Z����^��֒p�T��&2)�drw`�v��RUw��/���U�v�'6G��/�w`��b~�*sC�A�������)��d��d�
�~(�;*GLj�=�OR!ޗP�:xx�&P@ïq+s�D0!J�1���z�r�eȉ��<jQ l����p��NAd�m�j�L���ߠ�A�pG��x][>`�ί�_����[B���^�Ji�;��t�FA��[of�\����fo����L�ۭ��U�8�;����b���Ԝ��{D��ej�[��NXj�]].Q�q���љYˌ�h��ƫA�ͳ��!�<D:�r����:��3:��	GiVY���ٰo�^$=3�Yp��P9�����XF|X��>:��؍��TΖ�����i��R�2����1��P���L���^�@z]��FCz���祷M����%n�0�	���my_P/b���RD/r��ߜ���cc4qk�zZ�z���'��Ig�!t|��WA]�M cjʹ�
IH�˾�f���A������4tz ��-��a I��oxpk�1�Br�f����K�7��{����������3��V�pbKY(;4�Z��-�S�����O�Qd������+��e�1��v�8E���#*�v&Z���X߁�V?�]�6CE UFR�i��ɥ��r8YN�c�Xz����������a�Dy`�k2��8� �c�%%%4�=�E����ك��r~f�'�R+���J���*�L����('��0�dwi���\"�BUud0K�B�CB�Ѻ,
b��"�6I���s?�Յ��F�Wם�ɦq7PH/�սD5���lPXm��!K܂�%��	����	'�o��pJ�ʂ�D�e?�ل�,֍�G��(�\�ݔ��=L�����K�ԕ���X"�=�NFhp^��=�/��yV��Z_n�zq@?�[I鐅���@]�<x�Z�^73�i�.�(�X��;�[i�>i���K���
�m���I\����q�s�<Au'����]O�M[8^���,��� nn<q�7p��R[��d{��*F���J�;9��Wm�e'�J��Fư�h�:��˷�-2��ija6�e�Y�U�r����� ��@�:f4t�ᗑ��!�/a�6������uV���׆:�swZ��m=��A�@Y�jid��I[�}���w��t;����ho���J��$��i���
�}�F��6wK%�?'�����k~���z����c�)G��UL]Ub�&�""��@`�;� i�eP�|IO*w�����_ة4�g�n�����s����dLϾ|[���C�])
LX~`�7��q��_�>�C�=l�����6�"��`�$����%���VԀZԣB��_+���Te���l���'v@gRţ~���/�R�S�&� ՠ/D�GS�gJ:	�p/��H�F�o���P@���?\�TBz˛�|~o!N�2���>��I�������l�m �F�������'Z��)4�`�[08_�";�O*9�L6Y��;B@;)�G`�v���8���W39�,�2�5�UGL�j�~�zY���M�я}f]N1�'D{��}(k�&?��#�uuq��$#�)�i���<�]ə(�o�_L&����^VC�_�|W��a\���#9����J�g{D���%��7����`^tpab�ֈ�,��?�"<�<8�ƾO�Jk������0d�TK�Y�n˻�Y_	U`p�a�$5��le��nX^��:�>�S��Ol��ϝ�/{iUt��D:��=aZ����M�iY�鬝�;��g����2ѫ�r�AA�cY�pȘ�5��+�Zdc���@Т��4�͗<������zr���-�I�-���ｇ,����U@��&�|#��FՃ�	�c��֣3e�GQ��հ}���F+ANr����,T�Vm%K�:�L���eio�#v�lq���T�L>aK4��|#�O@�������� Jm�}�OO���v:g4t�I�U=�6?��O�l��)i%daP��:&WׁλTvƺ)��L���������b��!q�s������1*�P+F��X�O�(L���Zi���(/>J)ѱ=��v�Ā������:_�P4_E���B[(�nDN�3�StA�r�J��,oX��n�f���옫���Nt�&N��j�ˁ��x�M��C{���� t�N�r�j��g��ez����7_2=�h�h����\qܘ)o�q�`l`Ӵ�{����I2����+����wh����#�H� P>'b�A�d�3v+�A��U������b%f����L�R0[�whN��� s$�ϸ��x����cK]z �;n�Lm���v
��'ՋHӔ�V$)�P��揬�D�"�/��P9Z6Uvf�k�j��K��7���3��_ۨ��C$�7����=�YĒ�������yo=~Ʋ�Qv��?�)r��	� ��3I��^H��L��%�ν�B���fP��"����VB�JBz͙]!�<~��� }zR�Z?ɺx�z2�攫�⎃�w8h��@���W�E}e����l^�'�A��f{�]�`��6�Z�� �c��q�UR�o-^W���������6������t�G��{��16,މt�Q��O��a'e"q��V��Jy+�:��p;���w��P��;��YW�h(��?Kq��`7�
F{�6�#E@/O?*u��D�>�8xDQѲt*�T�������(I�Ĥp`F�:C�.D���F}z<������srJl��N��9�M0{��?d�����d<��Dݢ.�52���j�_w)�W�!9B�C�6�I�X'���5j�2�9#���&��[I�+��~[&���҉�(7e&K�c�U�uG��=��X\�pH<�5'�~�҇�5
v�`[6@h�(���n�s�|�4QV���K�J�����¹����"����\�v�	�h��X(��)��,�{	�LQL�!�l0��f��:���A@�i�3��xr,~	^�vd�-�:_�<�Dd��#K!1�{t����Rn�n����;���)������-��S�7�����S�X���}�۳<E�<��_I����5b���eMp�4x��'Zs��>����$d$��睤��!=��`�����8ʻ��t����y%L���@��k�Sf���f�u�wc�q]���ɓ]\'�l�B� �/b�w�Iڜ���A ���HW�d�E�k�/��%՞����әh�7`lj"'ߓ^婄�h(�S��yz$@���Cj ���	X�C�Q� �s7A&��8�Τ� M���w�6��]�MnyRR�t?�a����V�g���+���4����z2�H���#��g�J6&L��JX�ㄷ�V�Q_]:o<a�����h���C�Z��t������l(�$1���2��eR�R����D�^���\��ƐB�t�VIz�R���R�$H0��t[�z�Q��Bw���Yuf&��;����8�&|�#;�v��ޑ��x�3�Z���w�����Ex�%ѿsK��#�9�vZ�?�����:X�9I*⧯
)��?�G5d�˒��d5�_S�!�L�����]��r��)P%BOz��e�?��)�$�R����C!~Ͱ��<���Ƅ���Qs"�r/�7�G�&�/�)�x3�o{3v�7��wF�N�%�F�^�g.��br��� ���_�A�cC�����%�}�E[����W�Ç�k�G�����|J�^h�^�e	X��Ɇ}�A���������4���\��f���lD��/�����yK�1BكW��❾𮣨�Q�X!RF���oVT@�,�����c<�k�׸0���/�ZO�&���ۉ~�]ä�����eJ6/
4�� ظV.��K�N\4�������*��!���Dt���T׏
�-� ��)zP�i�2�p���`�j��֫�y����4�_����V�C�\����wj�t��{��3Z�ղ'��P�P��pa�|�����N�k���I]U|��~���*��m��g;�?Vg�3s�\��8Fx�oŏ=��fwk�U��f@��^�H��mŊ2��/-�|�1}����n���#�-8���M�٠h�e�[�����p_�0�h ��*Q"в}�d��:6c�[i%�NT�3�ɫ�%�E���R�I�����a|��³κ	��L� �u�x����)K�S���+:7<���>������_�}xC�B\�_��G�O-�y�Zփ1��!�(���3An���� G�r�h���ϫ{�_y����:di����7������s	u�صn���I��F�B|�,���ND3��e���)��͆r��Q�+Ƃ�;Y�I=&�+[by��Ï�bvjw��i��G��������?^��9j9�q?���,RN�2/+����-�;x��������Fߢ��k�p�YA�[P����}~�"f�V2��b2}<���PIs��'�)|Z��a5�)te�~R�Ql�N�(�B=�`��(�v��&�:�Hr� �g��߸����c��eRM�I�U�I�zӍ���ι��A>U�-���sF�}��dΏ_[<͹ZO�x���ҫ(̃�F��W���/�f�~����k��J��s1�y�^r�~W��!�\��Zܗ���e5�I���Fܸ���=ֈ?��Ui��&�$J��v��Wl�MT�RL�܊�<��ҵΖ��+�<�,����0�Ȝ>�W�2&1]�{}t8��(~�Cx��C��0<�Q�T�9� ����lreQ�du���$�c��q~��g�"���Z��Z�����,���pά���>+�������ք��\�|��W�0�2��$k=�$9��9���t�]W%,%�7�˲�@��3䠝�Nr����nƮ!4P;�}ANE��L-����1�Z(l��k�V#l���~}����^[0\� *�I'K���c�X�hc���Ҋ�V����! ��������2�����.��s�\����+X��[�<��؝�s���k�[??^*��}O��z���D��W�Pk��t���>�Tp[r�}���3�2�p���Ո&	�K����[ 1�sc��؄
k�tג��fO�3��E3">=�i?9�'~y�b
������y0o�����o<J^���L��N��X_G�o�0�@�<4��j/�P�dO,�c��� 7]�&�~�5��H�\
�c �C4e��:Y���}@��H�1E���5���tK�1qnA=���v
6)�0F e�-̰�p����E'R��`H.o���w�>2��X��8���s��8�V���_�=��w���I����N�U��w�N�[��ǟ׫�/ԋ�|�Jz�H[&�[vrV3�CH�g=Li��^3)�Zղ�7Y01w5��ؑf;`�� ��%�{9{J��˿L>���f3
�>��g$�\���zǀ���P,�ʳ;�������>�V��$�^�FH�|�O*�H2�?�z�cx�>j��3���^�jA	��:���c�A� �!M5�����+�m�R��(�s�������/#ZLP�ɂ��y��
5)*�e�q�	��{�(2����R�5C�4�&�H���)Bxe���1|�O�� /!��[Ii��Pl�O?ɤ�K���0_;;��jA���؛�Kފ����^.�#&��ȴ�#��,�f��Lk`��1)�~	?%�z�� ����O1�['F��i���� �Z���Q���Hv�����XUE6;����S���HN-��}�BU����8��E+�����c���������n�\�Db�
���$�{����ʈ�Ѓ'�ج�o��U)E�I�0�2Im3��c a�h.T9��s6A�]7㲁����h3�Ao�����r=�>qu����[���/H]G��\�{�ٸ\�X\�P�OJ1�*JA;�C���82��!؝�=�G­JQ�V��PLR�ᱤAS��`�5�>�n�Ŏb�������޼�:j�ƕ�tŹv��	���Z����qj����H[�`kEv�����t$T�ٵîJE���]��~��N���i�����Q���|����1��n;v��Η/�#i�������q���S�;����;ꋕ/�
�_�5I�x����ܨ�.�P-\�̹
Y6ݎi+:4�T7��]f�U�T��N�7fC�!)������Hi�|A��,�6�_�+8ܚa�N���@��,^G���s��y���Z�u1�AZgc�V��eW ��g��t���Bl��F���o϶ǹ��j������M趒�f6�����/��۟����.�Z�~<�y���h�wJ��P`F�|s�kM��ϲׁF���elM�K:c���A������/c� ����>��c�Jr�K�s�rN(�W�zw�0�H%cj5z;�?�P��OP����.��X��aCi{f�H��%r��ճ� ��hhU�$�
�!�慁�g�J
:���T'&�|�#[�2�'%cV:ŧO��/�i���3��`X����J�+���6�J�����"T����-̸}\��Wm�|���g��zJ�{�4�������l�k��QRrc������T*O�3�UEEE[�� 
�����^��5�Јd\�R_�i%�c61D��QE&B���!�O���x�3!�W����I���qɿ��[� ��7��7Z����U��r�iڃ����;�ҩ2���г��㊆ZF�^�G�{�	A���<){"�D�����O.vx3�m��F��Ɠ�v�Q�z*�:��M��v��:fi]qd0��^֣��v;�y����.y�,4�O�@o{���Y�ʏɢ:�}w|(�d&q�KG�:�:������̘y-���c a�<n��%N�+���i��(+{`�5m���;|l�^�������u(��ncF�T�4j	�.���,��D'�Uh����[�ײk�/ ew2�(L��2?��^-�HH�ۉ,c5w�bʿ�����3oQ�� %�q�<!9|�	*��u9��l�k%�Kk>��xy���iH�IM�/�����*�D���OϽ�+�H�l����������9-���֣��%9�����v����;��4	�T�����Qx�X���'��?�[Ƥ��jjPWjJx�v��3��˸��|֓Jr�$�w�kť�(Y���P�y�nK0�3 �ٍpڣ���=��K �#1��G��տ�X]?��?T.Y?V���X
s��t{<�:5 Ī�[a��|�y=����[�xmJ��|�א�`�f䫰�롲�!EE�Pp
w�Y(�2~�@ ��@K��VZ-f���0�ލ �Rǘ%�)bQ���,�a���K�<9�E�y���h_���|AO�,�M��z�.�<M?~�P6��Y�_��B��{�n������0�ƃ�	D��c�� �F��ה6�^�D.8��cPy��"[�����#p%A�Od�Ƀw� K�y�BAS��{�s����9���;��p%��"����M�LҺ�z�Y���&�\���ZC:)Q�H�mU �f�@���8�qp�2���(tc���((tH�n�~�����ފ�5^�q ��M��!�W�p<]�X,�P j0�%p��i�X��4���+��f;�YU�]�K+-)!iTf���+�?7�
-q�,dtr�x�~A���� ��'������qk���އ<�a^<�u?,��q�ߦ׏���W��^�)�o�k��A��PU�=��mߩ�H����۲���-�)���0�,Q��)�{��<�w��Z�%�Ma� L�B'�n��di�<�e��y�<�e�^�Yno؃�u?l*���o��VWl��~���1��zP�Ys������p�x��s�%��S�:����֐�W	�m�^#{���b�MG
t�K�\���q9�f=_xp�lT	i��voF�@E2q�*8�� ��0������p�&_��1A�D����eK�J���ӟ_�Յ�yL��	Y�B�e��a}�ݯI���.�Q���M6���O��P:�f�d��u�Pd5e�جJ@ %��7N
.���}5�m2[�:����uC��ώ��U��gL|�oH��I�����?&!M�]��`�j�L2(e�>�v{�yxX%��S��m�������g��?�w��~nŊ���5J��֕�r�ͪ���K�n���]ש�����{=%�>^����D�&��p�V7^���矁 ���΀�ŜV1�=\5�����9��˺�{���$��b�*���d��j�h�	4ڊ1R�L�������^��#�-�jFs��V�e�|���#�;DY�o�9pr�p��'��&�{�%�|4���V����W��������j�q(���u�J����wj�v�#"l�ڙ�7@&a�
R�<�����}#���p��'hn6k��CEj�z�\���;�|���)/���H)z�[�GE���T�Q�]���겲9y��V[�
�#��:M�&��C0O�>�*w#ֻq�b-�đ��]ok�?�P�gϔu�b�`��'F�?�N�w�AϞ��>�:)�A��V���CC��~�aǇ�aJ����@i;w��d����~R��Ճ��#��({3�h'FxU�`V�Y������S�����~��ek%2x(!�͓!�ypBP��0=�
�;�m #�ZW^���^�3�j*�G�*c,f,/O�p�@���(Φ���m39���Q�G��j�t��;�zC��Љ#y�5���r���Ʋn�N����*~��6.~m0�F��/o{^1AЇ��X�c�.=�:���vZ �)�pK������Xy3��켴���ׯ_M��ތlY�8�X�2���.{�82o09r�:���!KBLcc|��&�#@?���E�)�j��PZִ2��j�<� C��9�_�(/~v ��
5�g
���h���=���R)%�U�{��h�65c��l��Q���U@}H4	�|B�VZE�����S��T欢�"��)����	���ॖ�v|r\|%�z���#�/�	�_�h~{8��ה����R�Bk��H���[���H5��RbD��גB{p�$�*���k	4�N떇���ݦ���������H4�(�C�
#4�~Ȓ\�FV�]�̭@�G/[�?&2Et �ӷ�f��jA�+=����Ͼ������N�+^�#U�^U���/PHP����+Z�^]warsd	�φ[�4�74��5w��+����ePY��u�����Q��'�Ɂ�wˈ�h�����T���W!���i�+�$�I�{Al YMlt��o=��ڎ�C��ё�4��9��o���=��c��/|����~�ЋL(��bԕV5�:�S`���|�����{e��o�w�K�e�z�D��^?� ,�O�=�Z����R��|.%�G���VFܗպ��p�)�˨�K!�gIHd������R�y���֚����C�� ��ן�B�+�?z����t/���	B�`��GA�� �A�@�q��~��E���]FAX���5l7�����3���������������Rf���K'�v6��4��:�i͈�#��d[�W%�Z�c�':���G����FG�EӰf�"�3�盶>�3<u��>C��僡?��p �~�Z;,�����L�	?�蕱�ezD��X����U�P@zB������Snr����J���㷴����o0�!���U10�)���Қ@�C�Q�e��S��*��ȮoLtc�We��7�Ņ��9\��_��Xi�����������ï�=D��^�q[�v���ѷ���.38ʉ�1���Y�J�V�n���7=jXrrOFU�r��l��W���ܭQ{����uK�O��Μ�s�v�N�_%l�!E�����|�_V[�KƳ�Ijd�o&,S����=�����H�	�\�I���z��Z����wH���_��k�I�k�/
Lҝed�֝t
����I���-�^�hmG���IKGް��+O�؏�d��l ��"�~7ɯnF�����ͣ2oA��$4�{��[�Ib	i�$� s��Ϸä�7��U���bR���7If����++���f��df�8�;��S�"��eR̬\B97;i��>����n26�U%au���q"��B(��gIR�B<��pj��
�p��O����hζN��WU:�'�ꛙp�� �zK#���!��P��-�k�v�ۣ��ƛ@_G~��=�������6�[@��m����G�i!�k��Ү����/"���Q�P�pmy&CiQ�Ƀ#�d��~����L!���`��+L�A�ji�8�ݓ� -����唥���מB��4-?��a�8��s�#v��3�&��ŋ��E�%[���i0�#��T1�i�z��5&ɗsc�mw��=o�(ռ~� =�oX�5�\��C/�1���a�����s}�+���1?j_<ޚ��u���^���64�D� ��ń�s)��80�)ג �\��7F�����H)V(ӈά�����4��H5���y�φQ���e��]��;+�;�bX�E)|H��')jڊ6�d���9�C�Vp����:�%L��8��H����Ԗ�O�ev�����g61!Z/�l �bOŸ�n�Kgʓ]�Rn#�@Bi���%P$c^��%�q���:.���բ�XH
�^MZ]��}�(D°�k:1�[]������=�r#?�09�
*�;�G#0�j��T?ت����Q�d���m�G6���5�q��i���u��T	���g�`'�!�צ�.��
񼌔$��Pb�.�������"x/Ue̔@JHC�o�k�?3f!�c� G+|���Ɨ��nߦ�@���.AD��چwޛޓNC�~Ս"�GS}
�D��Hț)K�K���3*}�j���vh�8/`�J@�ދ4'���p�?����R_q��.	�8�XtBf�ϒ����yn�t��Ɉ�j�rn�vu��d���V@�4�n-�o.�eXXx��CšTF+KJ�Կr���\�3�%�b��P����FG�F��f��"�"��*c�U�3��>殐,G�����	Nf����T4��M��G��Fem�4٤�爊a�=���ഞ��bsg�#���P�#�#��d�vTy���3��%�Z%�:�޾���%5-&��Sg���p�X�`#'��G�xz�7*��2q�r����o���=��h��>킷��М���>Xv-������{�͞ܥ�Z�{��ko�{HgU����X�}t�R��7�O�}���ߌ��k�D��3#0�D��SA�]I��]-YIG� m`rץ�9�"���ߚ�8X#X-�=`i�d,Q�M���Ua�S7���j��1�Ǝu��&-�P���Ʋ�D�����!E�b���{$�1��=D�Ыn�ju���',*��
絶#��������u*��Դ��i����d��amj��y�/�r�X�^ߎ�wri��o*X�:��=�e�qΝZO�|�c��K�ED��-�䟅��"�S�H�w#�Q��+qCg�@({�7I%R4�r�ア�#N���u$7U�h!K�׳�T!hŧ�UMa�A/�,ozt����1ܦ���L"���%p����G�cG����b�l��\��-��Yx9R�Mt��~j ���VV�@�����Z!V���������{C�o��ه|=	8z���:U�?����	�Ln��h��f%Z�=�+�c��|����T��� :H�=�p#�u>*<�7Y��tձV��[@���O9����s�?nn��T����`����t�x
(b���`:!M���q�[�riD1\(��>��yH��A!�[�p�p,����#��%�Et{�q�1��ܿ�O_�d۾M���6��VAb��A�Q*��`0�K$DJ-Hw��*-"!%����}��_�y]��y\��|�	.ѳ�����3�7�d�v7$�ФIF3<�o��]n��&��9�W�?��䧪�+�0l���u:���YǟI/�g]`KN��J��p����c_��9���[;��]*~���8���r�H��j��X�
���3x�`0�������gw�\��I��f=�n��r/����9��EL�,v�@sF���a�vz�M�dl��#V�����Ѣ�s%��+�V�?J��e���~�@SHKB�R����8�D��P��������#В����Z9˙ݳ�-D���,��L�n*��������Zmh=:�f�V7�t}������/���-�E���mȫ��<�~-��.�1���v��q�{���Y
~�Nr3}�]�_��拽�����%�3���B�o������c�������DiD�=��Fc���,�d�Wc�zhGC����_��]�KS��.8T�ʏp^�F<����������0n=�GN3U�^��=����F�[�M�`5��l�;M��|4*?3��9�mk"@I�
�`�p�iY���nW�GL��m��ޗں�r�Ĥ���[y��b!��_�L�ٷ��4+��ow��N���a��j<����4Y�;Yo��c�����%���&���}�A��s,w�'��gHb�p}����>� Ѧ� =$�s���eԦD�,�QO���_��"��̒�(v?T�Z�L�JQ��4i��Ïb���m��d�yO@�F<�[�C����	]�_�T���P]hJU��R75/���4���$���늬�ڡW�~�u��9Ϝ��K�vh3C�Z����c��aWw���Iؼ������ME��yϹ/Ui�C��?Mk�y����}ϒr���v���=�Ւ���5��Ɔ�����5xwu~���)/�o4ǻ��f��$Q��В���d�x�(|ZT�a�cU���z��(j�G�E�,�k���))j�p�6 �%<�r��L���k�m]5j���h
{�)��0,�5O��y�h�U�S�;I��K���c�?m����:�����2��!����Q������.��=�b��𹏀|b��x3�+=��)�M��!@	ZPos��*H�g��շ�]��RG�ѷ���ʥ�D{�K�:F5xmX���!����L+�) �N�3�b3�Z΁q�c_���ӈ����k�	�ĊD�Έ}8Dw���8�O�ԑ�{�Y�;��W�I[�-S�G��F��0��\�|�"Ie8䬃Dc-�R�$N�v><vU���ۑD�����l��:��8�9���XU�G��a�8��?����(���
j�OEz�m7�[�@���2Six������|RV#�ve@�y򲛾���{s4�A�\6g�ߴ��G~��D���PR�N���r�^�����r
��W����X�:U�Y������1�������?m$C&����.���;C�h]��T�"�=(�<������?��^SAp��<}"�Z4��0Ц&n���W�ӶEn��A����Q>?_�:�]tHOU���$2s�,5>�"�]
�$w�ڮS��߿Z7��rx�c����;���0nBK������x@{��AL����Ί�LV�9�c���]o}*\%���o&��*,k��#���@J�6 %u .E�n��4n)���t�tŀ7b�����i���ċo�I�
Pv"��7�Y�&���)z���e��&���6Z�������g]%V���9)הW���T�7L	�һٺ�*�~�4���wW�E�U��%*lż�ʟL!(�Q_:_����{]8�h�G�C3������T��%_%��������'��$�у�N��+�|���n�Nwf�sAw*w%����qf3���M$I�:�))��������]�>�$�)�N��QU�m��� IZ+}�\v���~Z�=�鮘l+��pF�W! ����R�T���t�>v�z� 9I��X�'���/8�E>�2?�U��=р�]�5�w6:���)���q���������:��_��/�(��Q��������p��P��k؃8Ħ^s�!}Tw�~g�qC��&l��/g�ӫI���8�
���j����5��o�9���p�/��A@�~���:ڿs2�8+�u�0��$5Q��ׇ�#[�[,ܤ}6���v��{�0C�����rB�JH�˥�OAH��\�7�5��X�ZE�PG��=�?��>1*9��m����!M�,�	3t��F6�s�E�������ۇ���nyT$Еu�<���a�gd.آN�,�5���q�%*��@{+��m�Yoz�5��ο�����
�
?������������6N�,�4��Wev�M�W[�"^�^Ld9���t:�ݦg'Mr������B.
<��
�����K�x?���̼��Z]ߙXW�Ad�C��*����}=��N^w	�+��!@'����f?۪(��"\B�V������;��V���8���d�@~��j�]�� �%��} �l���s5�,��wf�(+��k6n6r��)�u]ߚ�u�hBA�ةP "�����-��
~{�	����m)�ݻ�,��v���`��
�9`d#�,�|���7��f�ph���<쭬��Go�x�P����@CB����=L>�*�!�B��a����'�z�v\���:"��,�g�a<Y�F�t����?>�c�ͧ?����ڶ����l�1翙�\�w���ct �������UC�k+�A��3�Y4�5�G�7�L\E�P��L��"�����n$r쨯��$�\�Tޡ�Lq�cާ�Fq�aH��..Y����e��)���Ͽ����Ӑٲ��,�o��F�qn=�]l4<�T�Mk�X}@K<������~�:���4��~:�o�B����Z��@�W/�N61�$L��Ĉ��Do�/&��e1�9�(	��F�>ńX�A�֬�z��L�'�ۓ1E����� ��9��f�<��T;&�ХԂ����t����ZwhV��� �-y�U)��`��?�<a��`nQ�'4���qoB��e����X?.n�����ea��?��V�Smv�}����R����ڥM�6�`y�|c;}5�FQ��	t� ��$�wc�W��ƃs3q�ײ|��l�_�,<vxܠ�D4oѼ�vʏ������� �8]����gHl��X���p�)R�1Q?�.�7�%
��o(��������b�)3Ƕ;��[�uuν�"����?'������S�B��
I��e���x�i������@枾���)�d�a�F�Li%����":�~"��&�9�[�/(9{�I�g��>ݺ-^q�b�V}Xk�f����tɲ��9�N��Bư���Ǽ� Q�&���s>���"�_.T"�v�@uHt��D6���3
S�#���(� s_<D�*�Äd�[7���-�݄O�|5���b�*|b||�����OЯ��J��vkgL�*N���U��J��V�����Nq�P�.�r���ÕV*i^C&
�X��ҧ�`�9��W��?E��>����E�?֢��m"�#�6���
���K��8œ��R��A'�~���x���NB��v�����U����RjcG���H"B��tg^��"�����Y �$u9����|~���Ԁ ���X��������,^��VMu�p�-�S�&ߡ��v�VƱ~�����zx�~3|;���W��0�e[����#��q*
yDśͮ�!�ӭ�R�v|+�Q��B=��� �zL�H�Ռ����B��-x�0)��O�wa{�Nu�E�I��	Ͷ_|���ْ�'�����%���LA0�ȯ��D;5ڧo���vMN�Ni�3&R�\vt<t\�}ϊ��,q�#3l�����t,2)��r���v�<j��*hH��r���qTUK�c�HT�~�������z��Z�#q���/�Đ���9� W�|� 5�??�C�h����߾��ayD�v��o�w9oJ��4	��${G+ޚ��v�,/�E�Iڣ���e��X��$>�z3|c8���]w���{���7�m�#���~���
$�K���F�������5���T76c&.i����b��Ƃ�S4���ƒ�v��F$ƖɨOn�0�h�� �"^���6��t:���V�f�'+m����f0�ˀ����V�?ʀ�y��y,+�lW_3[7W?���~���OB��_8%r�[M'2�J��Z<پ�t
�`a����a`G�-ޠ����Ax���|�I��w��I����{xd6�N6&�$�A4M,ES�g�A�@IM)պ��Έ hEX�������Af�wY�~邗��,�B�PJ�q��ɐ$�s6Ů�,Hɇp��;I�p#�_�U�'Wb,��٥��L[;i�X=(��n��ʜwG-�ȟ��s܎`w h�$�ِl@J��y��[3���t{�N���������J9��g�s��Fj�B߻��u]�8*g�X�uCKT�9_Q7�І������i��C�ҡ	g&��{�D����w9~_��� ڜP�QB�-94��E4����W��݉U��ӕ�;Η�Z�`�P����ՌF޿ Z�l� �hQ 1���#�jh�rlV9M@��������oQ�����	��~t�o_�.�LF���S�Ii 6�(E��YM{�)��<���-��V����0���2�#D;n�b(Pj0f�/�(ЂY~�)��~���±r�q���, 7���.ܝ%k���F�O�(^��:b��^zd��[�'�Kp�5L����j(�\�4�z3GƬ3dg��>k��J(�0f�88�Ţn�DD�3���O'�2Ύł���SL��pb�����8S%�[� ^�a4�'�ﵶ�����S奯*IK��;�9��ǋ>�.]��[�C�I�>���P�:�E�Z5�I��Ḥ7L�!%S�"Nf�Cupѝ���]���x��U�}���\ُ5�W��%���9��$�n�HE���d����Y��Q���%�~0���C�$�����^��'���o�����kȢŖ���|N���I��`���c�]���Tb�|Tn0R��,�`�#�[�Ϸ����IHX��񻟵��S�7��-���,��� ��o)�+���zL�@�B��|Е{�%1�W@�8�,�]�c����#R�y<�>zU��ӥ��:hy`:����H�0��5�s�UU�<�fgaL���S��7o?K�|��宫�d]��7�1��	M�҂�V���!��G��5��>���q۟���{��fl&���m]^z��zH�.y�}/��=.��7h/6K�Vf+�s�&R�j�� na�uZa���:~/6z�4!CN��3pi�.�x��x[����x�&�! �G�Fs�߱cO�T�>�#�Da+\Œ�jR���w�
�Iǚ�Q��K�x�Q��Հ��v���F	~��%��Om�^Yj�jͥ�2��/R�.rH�4�T��D��I���'��p=��j�1}��p1-���PR;x����DW�
�����x��/���$u�TnKFn�2��g�b�x}����p����g8��<�op�hv͛���y����V
��4�g[S���/��� 8���`��?[���;8��^AW��V���W�G���?��r��^+�o�jp�'B?\��PͮD%ȧ�L�j<����)i�T�"t�P~�Lf|&@3�㥋z�nQ{��,Sڧ�`hiӫs�C�[�D5��fu�)#EO�QZ�[jċĀ5Tl���B����f]���Us�Jћp*͙ݕ|�4����'�k�ju���R��Dx����t�)��t��;n��XR���c�׶<�n\�V�M���� �l��;}�V�[ٍ?p#�����`��_�dV[�w����7�}�;C?�?S�����}�����D��y.�}%L�&��S�]���qݯe}'l5X��u������xoJO��92*�iHB��#s(U[i�(
�����r�(�tكy�h��v fD��i5bN��C>���uB���Ră��Ù�c�������!��O��8RVAC�U�=~�é��(LD""�%��$]��럶*t7�/o�8�J￥���:"��=����	�����R�����g+
��V��W>�R�r�KrUi�)OK_T�n�F�e�8��,���2�8X ֯�C"��W�NM?�z����p~|��w���x�˖?Y�����w��$�%�_Jo��մ���-���9u����'�
��(���w�5�1��6Zt@.,�������vkB��G�J��
��t�,��	)ܳ.hY�	�<d=1 ��ɯS��8ra�Vxޕ�HTJ�$L?�]��*xC)�m��Ij�&�v t��D�l�,�Sx?�l�ݓ��Z��>uR�b��h���o��e �E�>����i�Q���5N�՞*���dMU��/�&V���5���E8�c+Z#@����(}ЩZ�{���c��ZvGff�SIK�����h�@�u`���ͫ�w�ǲ�>����9T���~���-j�����.o�/������*�;���~q.t���L�Aw$��tD��2и٨6!�|#V�����|uH�jD�F�B�}#�|F�"��$�h�L�OU��I5�gx\��T��A����b��"z�V"V$ۡ����-���vV��ǋ�^�l�$�����J�"ɽ��l�|p&R'�:�v<<}'.�Օ�8h��EpU���f0�i�}���dN�hdm����$�W{��d����h���/�o��KuY�g��
���>�S��8������A��X���]/�j1~N��Rx� Z��z��ź��E�b��.�/�<��5�yAFRr�۶X��h{�Y-ˎ������ ϫ�\^��G�2١�c���v+��D��ǎ}�^��{x5��"������5/_�����U�s���cC����03AR��z���c����&����nKOg��)@}�����Uaz�Ȝ�	�'$,&o��X���$\,�a(��^�^ٳ]���p�d���E}g� �GܧS��c׾��tF�˧�~h�����1Jb8��3tM�UEmAE�ˡ
	�T:�Nj�M=�a8�r�q�M���#�'rM����o���^H�f�s�U}���>��)d��7Z��v'�=P�`W0H�{v���U���y^C�rWÁ��=�Ț���,1g�ؚ���o-+�3U��aiU��%��Ǒ:H�>�#����X���L����}6��n��ӧy2{������d���/�W��Y�~F];��ʑ���˶.^��x��v/ ^�k�Y<c8[����߅��3Δ���u��~kxO��"OID��PV LQ���k����f���{Mk"X�oY�I^��*h��`�bC�W _��f
JXgn@���"6�
��Fr9�Fv��Q�RG��o�|w�� �ۼk�0�*�.y���h�"���h*X�4���E�=�Z�f^m��XL��w��F�e�H-� A�#�k���)���#2�q�m�Sg ��X�vC��,��N�yZ�
S�۸�����_�8�>�5�����c�<2&u/�t�f��	6�B��P`�F&m��[G��u٦�)�W?�D�h��mot��w������t/x<W7t��v>���_61��ONNKO��|8C<Ǚaap_�?݋9�����+������_^ng ���PdNҵa���a�)*�t���fe���q�)�Ô�U�h�èf�>4��fI�g���n����1w"r�)"8�t���]���=�B�ԏ������������5���D��_Ff�#��(���줳�
t�A��SQ+�9!��I�����	{sw�Q���]/��^�K��T��S���m�Y��v���$Rߟ�
,�`3Z�$i��j>��]������'[zy�~�a8amǬ���&'����A�Ŵ2�jC�>*q�T�g��$� j-��R;%��H(U#N�棆YM�'s[�S������_LUe%g^�r�(�y8nث܌����\��C��~�<���˔����������ڡ�.��jc;��j�����F�e�?2��>�����q���&%N�3Xv��P	ܹp���}���%�[_���QWM�T��;��a�a�����^Y��~���/A�"����K��w�U��_@cFw��4�0��8}����U�fOu;�`8#��~`���nM�j"�y~}zu����b'�:�Ĩ���rnSM�NU=�u�c���c ����;bЦK}s���6���I�G��0w�R��o������8�>Z�(��!k�A�eAh��Z�����H���߲x(Ĳ����f�|���à���]�"1� �%�J�pKT�l�Ldf����U����\�}E�軹�.�j���g���󮬬���9�w��Zv�6�<e��I�w�7ǿ�ܷ��f��B-�	����J�����gn=������Z�:�'��f�x��j�f_\a��u���%�{R��M�ӀM�����4�6b�QC�u�z5�e��rd�[{~:J��#ɵ�����y�#�%Y�ư�%�<;�	��R��S
�(�X��rj����N��~---��_�7;ZB�m�ۣ�,�gB�=��1��87G��{��Mɋ����Tx�\�+WC�v��:)q̡L�:��%P���1��!�ݩ���/�Zh�����������!��;�p���t���OOq��R~y	S-��e\(�?���͐R�lu��<�����ƭ%2O�,~>Ҩ��n�~a���i���e�Up�o�0-��v�/�6Wޟ9����!�������G�dhUZ�nl�Ý�dtUa���A(�N�?#�$�U��IME���I��W4Tgtb�DHJ,�E�Z`E�o�1���� i�h��t�-}v�,��1�i�}��A�T�E�C���I�N��,|j𘓩�an��&��E�)�.	u"m9V(��\�1�����(�ij^"��BD�d���-(���ٗ�ՠ�>��`�����~ ����H���c/�	���s8�����и��w׳o��ց
a�x@�����l�3�7�A���@〖㩹�:�l#S��F	�3_ؽTx����qmT�����}ר֭'�!������=y��ػ�,���ףc���R����I-ɀ����;�'j��sY�p�r��=�#!	�qa!3�PdHd��a��;#oy�-
/VE��8��jg�����aI��G[�[Ҫ{T��4;�j>��}��jtZ>]�gJebq9D(d<ɮ�ux�H����KI�j��2��P�,ʥ�r6�#���@��*.�&���k2��<#�p�z��;��6��]<O�-�c��x0��n����~�L������O�iU"�v ��c9O}�)e�i��$�9&��Ѝs�~§Gh�nI%^�8]$A��\O9;�4���S�tӲ�3́k�^���0*M8�Ѳ3'����Н��/��3%ד��*�ʞ��<��&�_������pë�|'�g��9��V��筧<���m����Bz6+=>eI�IG�@
_Ai*)��",���ÌVc��E��)�����ZYT>u�H�ς�m�*�������<5X��ȸ�8��X:1�SCUR�9$�-�<��#v*m�rb��=B����WO�'������f�Ǒ�98j�G�"Ζ9�� �o�5��#&U��L�Pr��=���&#�~xY��\�yh�u�|�N������*�wg�jLz�ΰ� ;���fpE�-u�T߮1v=�X���Л뻷����6��ʬ�*�"!�ɽ�L���w�1�w?`.�W%��)q%��B���Yļ�gG���E��!�<���G(�������}�w7Ҝ�.Nr��a:Y�启i�ֽ��4�W��߿�k�G�����,�~Tna�6g�udֲ�O�Ig� v[�F���M���mEbk�D�Q�6+j:D����k��m�5���P��|H��S������R����-�x-k�ҭ�.]g3տ)}������!�����<"ꂪՋ�E���`(Iؔ���pXk}-�%"��:`�@�v��;��a��j�p��I���A��Щ�k�i<���	8��lSAV6
_��8*�D]��e�^Z�鹦��質n������cw����O=���W �U|������>�Sy��D��jy\̊v7s_�J���6���E�iH�WC�����H���R�J��S������#�k���H�����w0��j��5=SK,���c�Bw��������ث0jG���	O�Ƹ�T����[ʘ�"���U���(B�5��D����{��?{_G��ع��K\%��V�Ķ�}3t/M+�ͼ�1���,���S�8Us�c�c����*�
�R�Wb%��dyC�?�����pi�r�(������|!@�ȨA��]��8���3�yﳾ��6�V��1�/� ��W$}5�FʙHϽE�f�m/9�h|�a�M�[��~���07���o`0�����ø?����A6w2N�z{h/å�[��\����>���}}05?O�s!��4=JN;�l�p�1?Q^Ꜫ���K~�0�'Z��ss���Ik>�eE$�լ(�U��ܒZ��F��t0�R���c��&��{+K<��z
/(ȥ��JT�9j�PL������p)K��%�F
�R��������T6\J���[�c9��i��_D�ψ����C&�(�y<����l(%�Y�}L��QJ�y�j{�I��`��X��MvG}�$�^?���J ����(HazT�ѷNA�@���mi��L:������ٓ��>�ـ|m�X|����퓿�C�����Wԟ�w���hH?b�q�<nu{�F4�1ߣRkٲ�v��=a,��|�]`W˲}�E@L�`k���.Y�$�{/~�
ԝ�-��q(M�}vf&�)H�����^M?�޻{� -O�h!G\�ܸ���nly+���e �6����c ����N�5�Zax�20n1�x��vW�K�)� o0��F-��.��Oڬ7�z:�UZ�B�;t��-X�Jr��P�\��$K�A?��?��쓥�g,����O����x\�h�CE���C��g���YO�H݁;O=hB=�,=�b�_V;��tK�ձ�NmG�7�W�I�F��j�$~��1M$���������A/[���E�`Y��U,H������iu�<��Y�I��<�gU�GV�~^!"����&��e�U�x&��$������U��u��J!���څ����1�&\�'Փ�?��;+���=x�>S�/(���P=��_�Vu#X��:Ӛ�������P������!}���[��,]�\*�����{�٧����{��"QXl���S&�Rm���q�����kd{[Dx��L�D�K#K1;+���#�r��\��q��F�.�cݛjK��t���E���� GN��S]�GlMܝ���x��{H�V����H����Nq����oX�C�d�H����J��e�誺��J�O���_l�����+-3��n�������{�!���#�:I	��w3���.�*���0 ��Z�ħ�56���^����p�Y�x�����DB���_Ȇ�����\0����厰��.��'1)?�\�I��|�˗W#�y�mWc��C�Y�m���E�* a0TXA� \���h28��i5�O͆ه"� ~Ko a�e���Nk
���)���N\�����R#��y#����ǘX�Y6���@h|9�������6\�.�pS*f���. r9*=�(Ԃ�w(�KgrX��W�8H�N�y��/c�! ��N�e�����dW�T��qV�-c)԰)����-{�i�5����������c�^�0�0ůg78�Jedck��ߴ<���h%�O���G���/�����Rț�����'ȻGY���Ō�,�d��#��Fu~G������ݑ�M��m�n�H:Ϥ���Z巊>��S�	�*R`y������i�E�QLt�\�0X@�B�ۚP]4���~#�����h�U`���6u�=7�����)!��S���2���+�"_�K�z#��ny���<�aQLv�����������%�zuW�w���f��auY���v7m�R�Sk"E/�� ��X���)�*jDl5��@49ΗrZg���\�//���}������Lwl�T��jIN7��B�XC������Bzo��U?�c��Ο*�up���W{c�%�*�}�ԃ{�[n�T��I2��<���e�
9
�B� ��d��v+b޷h�����1hUћ*`���bkJ�2,A>p�s�<Ǣ�eӴ�5QSUU�H5fljj:��KHU�Ɩ��p��jr:4x�
`U�} ��`
^�9 ��˺�x�JO�'ik�[���Ek�m�*OȘ�	_i�5���`'+G�C6���E�l^|	�h���?��P���n�Z,u,�/]��H0��L��Z��oV)u|1�!,i�Ks��<�����h+�k�uе���TH>�����Q�`n�1�`�qTV1\�����������]�5���"�$s��1|��lH��(��_%��m_���3[6rd*�T��=��z���%��{F䃣��\�W�Q��?}ײ�E�z����b҈:�,{;ՠ����d���v�;.�w���Q�i����]��/��'��}���VR��~���!�0�* {��������zD-J�&�͂Jj�k2՝��N&�M�^D�<'�>Z=�v?�%��AE�+H����W�޽,f���$����Ǭ����&�3$a��N9I@[��:��z>i��~o:ρ�}��E�{��^��T�P*�ܝ��f���6
���d�:q+q\}�����H���$u��}V�s�1~�'N� f}܇���t@�^��t�����C)�/t��>[���1?rz���c��=�����!���_�G��D�)�_�n��j��Lg�Cq��,M1�<���eM
�f���ߛ��7mrS��X��������;�+:�n���zz��;	�U����g {G� � ��%�з�f�>�6N��|�g�1D��rY�=�Ox��_-J�f|2n�d�`U��,9AW�m�ɢ8֞A���y�:��$�R�M9iw�u��y��tiӹb��{�UW�R�R�T�ݧ�@<Zvid������
��JA�=u���Y�|������\�gq�x֜��H�Z�3���`*^ڹ!W֪��z<��$�\Y�y�]�}�bC/S��>�\�ٲ���/9u�rTU�2�k�����H��K�V?��r�DW�<�DbH{�8�y���p�5�f���vg��$�o�^�Q$,=�G&m:C�R�G�@q�ތ���#X�F?�2vft��Ȓ3����\��可�pEhkWL(��Tg��mJ����ذ����y� ,��X��8�#��A�0�v߿�ͣp��-��K�|�R�	�T!Qi���������)�e��0�t�)��B#��L���iW��d�����$�_����5}�kq�}JK�?skz����8�KP�`"Vml�F�*̰�\8�T8[���쓆�@	5:���=�������+=ۙ�!�~�����U�ҕ[�~V�6��a�.����3%y	%y��F�TZ�L��I����f�}B��|SQ��#�����N�=gҗ��s���Ǜ�Qd4�r���J4��q����+�7����s��Z�
���=�ŗ�0��� V���5Z+j�t�y:��h����� �,��ƺ�ӿ��O��Q���ΝL�}��?�!��6B�d[k�f� Id7��T������	� 5����A��c/Ö�)�ڀ��fW#����ey'ML��[����s��U�w��8'��T�d�FuH�8�FZ�ox�yE�T�[��avS���pH��fR�0#�(_�F�yz�Z0[�s�KΟ71��s�9����<�?�)~��j�r����V����L��9i[aBmJ� W��9�K�9�7�H�Zrd���?��xN�k����{��y�V%$x�g���f����ؒ��(N��C�/$i��;��X���Ӽ
�	v��"[o��<9[���CV!(��QbX�c���F��'�f3ϫ3H�4�1S��o��P�K�Vh"VP7ZF�$M�fTvX�]B�L-�{�l�2q�2cb*� e�߉�I�_�*��6y8|US�3�2*uC@��{89V)x3`�=�ʁ|�4����8)�C1��Ř��9dJb�,V� �w�ڌ66�8���9���$��e�׫��lb����\��<s���
d��b��/lO�n���mJ4Pb�X~�ͱ��M��ϖ�G΅���:���ft��y�L����R��r4+ �!��J�׮M�����>�����J��z�^��	�Nte��!a�R�"K�E�rLDw�W%��z�jq�Wź��F]�ҡM��fI��<]1�!�t�T��S���J�P��3g�U��f���SN�u��WT���Ht�Yz��4N�Ĭ��eE�)�l�H����j�@��k�q9�C���}kB_/
�'��ʪk[�S�k�B��Qq$ˏ�����q<�Ǻ��L�&�})H�v9��g��>Ƚלw?��Z�3��}I�&Q!�,7��Y`ђ�|��������.���޶�������U�7%��m  ����:)�����t\�q����{�>}Z�%w*�q�������)gPw)�꒵�$�+mK��Y��'��	A��]@?Z	2;�NH���.C~�NQ���� `YV�����|�N��ڙI�Y�DLqs��Ž����$����l J6�Jڵ+i�A#���M氣Z�-QJ3�Cp�У�h�F�Vy!\;E[�����5:H�ݧ� ���.�E~5}�G�}i�J�ܧ��pg��9�)k�EE�
a�.�"n���x��&���lR�0!?�3�;�.�_o]��Ҳ2�>��E���cXdn|���>l{���6�͟��w�:��Թ��a��ӆ���sRI5j;��_��)E6�rI~�{}a���~x�*����`tZO���Ri��X��4�M���%2��|ff�^��bP0�I蛯���\�E�����6��PmfWJi (Z��p��:Q���M������3߮+Luܛ�5Kb�F�L�1��zg�]����5�x����`K�0u� ����k��/foEˌ�K�][�b2�s�3X��쐏��N�P�9<6�Z@���;>u.p]���@��2�R�N?>4���ϳ��|ij3HJt�1��K��Ċc�'��ej�v�x�)�8?m��ň=!F�m|����l�t��ycEy���LSs�v�q��:=�ũ�f���c����f3�X�He_�O��ҏ�!7W{��Ot����҃?��C�/+�_T:-}*�[s 2Ȯ�4�>X�?Q:����</g�����)H��NL�+��]⭜ҐѲ6��Я����\4w\zhR��סg�2-De2�KB�7 [b[Y��$t�j���K3�6��\q���h�� ����{���鈔f��7Q�@��=�b���`�i��s=s���R���o�)2�ú�����q��t��B�@�>��W������W50/�k���uC�nH�����ɥ��&�����g�����x��t���<7>3x���"qk�c���Oߍ�[i���ӥ���g�{�۟E�0�ǰW^I���Fsr�R��tM�W��?���j��zi�)e�x^���*K-ūf��v�Bd�ٓ��v�i��s��'4>�!�}s��8G	�ﯼs���"�OzY�H�����M]>zxqW-bj�ƚ]k����YOBmZ}#��X����@գ�e��]C�TvK�&a�'�ϒ"�:5+�5?�� ν+X�1����1_�ǩ����<#���+��8�U޿� ��fk��Zpq�q}�������w�QK��+�L���@�6V^=}�A;˛���\����+^_�N/���~�E}YXXh���|��%�ˡk\�O﯑Un�7E��xz�s�>_�j�dnU:o"\3��OCN2����|Y,hm��e��l�q����D}����B�����ڛ�K�ݴ��ݟ�0����LF��m]�[_,��?�qz�ߡ��23�&�*C�Jqj�n��1	���U�C����j 	݉E��и�T�!�����cҫ^�ҕF�JtTsV1�|��2��c��H�ҭi6w�'{���QuN�V%���x�k�&���y��TɊ�oLz��md����Q%t�S���qI���`�_�i]Bڌ�/��%�شΏp0Q7.!���y��½�T���A+�5u�@ ���l2��?��+��;�gi����x~�.��:���}}��w3/�YJ�{�-�U\�!c;*Y��ϴ�:��7*���,]{<���w�ӆ�]�r��/����}�r��EetS��ؐ�\"�ts��(w��[���*ʵ"�ｾ?�x�g��|�^���9��d���A������N�K��v#�ZLKK�pNN��|�{L�[�#L}���k>�nf��	�1��MRsy����B�q�C_�����3�|[�ɲ�#^�Z_��.�e�G��Ó��/L���{�=�T�	|��ic@�\&��{~l����p}&�847R��!����^B��ˀ�\��{;�j����Wǳ�Y�TA�ʓ
�Gټ
��=�~����<hC��o�Jrl4t�8����Gp�`0ɷ_��0�X�N�f�����^Jy�u�S��R��R;��{�!ۓt�����$���Zxfx��ާ'+���Ok|FZ���щ�=z�ݶX3ET��6|����?o�N*���D2D	~��n��[���4?�"�aN�z���KI�_+�|���mx{���wG>��K��;w���Z竤������Td
E�Bʟv�_�;�m�w��߫��*�{�MPj21���*��"*�`>J��k�I]ƃ��x=,��y4C�Kp���#Oxi�)ы5��K͔�\�B��Ev��JjJ)Bd�M�I�~��T�������A�.E���ˠݮ��U�� �?����qK�z�Ƚ�/��\�~�:G��Ę��z!��������d�{z��[��n�0��;␁��5�+;pt��|$gzq%ygs��L,��d\�����L����XP-��b4�o�8j�wo>���)U�p��+t���N������u���!����.��ㅧ.�[�������oy'�0\�����给��[7�ޱ����g�|������<�"w�5mB�O��\�����<��|8��?O]���$��p��F��W��CE��/�Գ*#"9W=[�..�0��
���2�b<���\t��sm��^���xҷ}�8���
�+�4���
�U1:g���+U���w���1���3}���A8���a7 q|��C-�$^���ӏ��.v�Rq�����+޳���{K���VA�(b5{�-O҅S5��m�g�- ~Ń�pA�� [�\��s����5kOݗ��:�B�x�_Z��X�Ѫٷ���;�%���]<�rpw����) �wc#ߟ���>vz�����f��������^�\(��]^,9�go��3TГ:$��␲�ƐQuv[���Qs��s�|גO��L��+�y��c�0i��ߒ��Q������/v�*E��@�~,x��&S>&�Z�?ty?�c���:��%#���T�T��}���RQ����&�;�o���ŕ��2��
x$��̊8�!�H��o�40F��q��BT��.�2A���(�r �x�׵�l�U}Hդ`b���]b�j�V]�̝��ۓ"���0���~=Oq����i�s�4@�
^�q��g���ƮQϝ�A)��WxI&�*+�HA���f���_�;����e5�X�����(<�q�]��~@u��c?2�<t��y؊8�~�e�RJDh{I)�,�+sy�,�*���ʲf~��5�'�[?�ܿ]f؟�/������fL�߀�[8�B�[���%��g�~��\4��o�x�!��sm��4���[��[��~[(���}ȇ�|�M>�H�����i]\�8O>U�s|n��):��C��'��G.��V�<I)b^��uv<�>Kk9����а�qr�(g��g7��j����s��G>��ϝ{���k>��������R�?��}��;d���p�L���RJu�h>y��k��O{�xJ� �G[���e�
R�K��\à����n]^e��3�pW����s_�9�}��P�Չᦢ�,�����A/2>�;��i)ڏx�H�ꢆ4
����f�W�T%&M7s��G���`�����q{b��!k`�����@��@fc�佀h�߇C�w����{/627Ȟ辤�ͧ��25�*������OÃُw��>6�
G�n�_�1[H��v�]�X*���t�/�U���CZF.M*���r���J���=j��o����O��jE��g@.\_��-kf�'��?���,����%�ŧ�H��'PjQK��ܮ�����}�Q§���P l��Z���o��0���J(1������o͓O�gD�gH74?�U[{T|�z���s�h���[����A}�zI����η��v[��J��~�c���ݔ_b��n^��k���[��l}<3Q��c�x�͔��V�)x^�go$]�c�3�ꃌ��#u-eHU��b��ɯ�F�m_:�k$��ld��8]d����8qh��d���\��?�
QF׭i�e�V�^$1A$9�I��;@�gO����\������\o���	j�D0�K����A��K	����ɵj<E� ��ׇ}�6������K�>�f$.�>�n���&Df���f�Ϛ_�s*	��r��J��߿C�j�Sj2\��~ys�qgG3����v�6k��������1l�������aܥ��C�u�Nw���4��պN�K�b=�p�lFj����=�8�����a�k�F�Ov��Ɛ����&E�.�ʌZ�>}�������?�������L|���%o����Υ���K%�:v�ϴ��~B?�g��{��Έ~��ӧ?��]��qx������i���#ж�.�P>�Oٻ���~nErOI%ߊ��~5�j�m� �}�ђ8ˊ�h�Jk8q]GbëG���J��Ёqz�Z"&3�u�_8�,˹�r'R+�s�\���\���Z�j� ��%��Œ�]�Z��<� �y
���i��[ kb�w������)3:�=��_X��Ƣ=��Ƶk8'���&Y�|���gi"�*¶D�<��MT�α��r��m�4$ً�����,��{�>)+a�|m����I��Mk���[�wN:�Υ���nÕ����Z}��w������wo�,�6��g�ץKcB��+�;��>��䗯�(<u���+Ŧ���+��ĥ�@�#Af��������s^<�'��W]�����_���}�د���Bf���/�9�`8��D|g����mj`�=�M�^��ѵ.��o�=R�~}��!N/��O�fq�ċ�w��'{�p� ���D��kfBƩ��&�5�"$�){���⠶�֤O�ɽOE�wf����%t��Z0�>�دف����0g��t���7���aq{q��R7���<]�֘|>q��І��f�|�ݬǕ��TX����͚W'��f�ɪ�J��4��j��ua�{�d"�/���v�L!�w-C�6�
�(��V���m��ę
�1���/V?�����:d�=��'U�L�4t�|t}���#;�̏��ʅ��| d������.�\c#��>����pvF4*WY��ʄ�<�c�z�����eWPJIw|7�|��
�aw�o�ɯZ�Cep��ߕҵ�}��vLwl�~���2�!|�p����I��6+]��������iUS�߃�K�e@��|����d��<R�|���iJ�G&%X�ws�lDA�{���M{�ϾƼ�?�StJ���J��o�9��X2o��l���{9�ِ��D��kS.&�~��se�Ƣ��!�&2� ��R��e�*w���J*��6G,�C�6��P��=k���2��qX��^ԏ9�G>���r)�w�3�pyO@�����Y=Կv�#���n�o�Q#�
�ZX���צ�Z�u-�4k������V[o��A��H�vƵ�.�?�IM_�z-����M�Y�z�2�	���|#�i�f�%FP��k�XZ^D���?�Q1"�zKƍ�kB;�����\>t���?�k[�.�(�7s��D{^Xl�����Ç��nY�V������N$�d�F�uw%\�{�Sb��"�g�Ti��(8�VU�5�1?;��FS�+�ktŃW֥��F����9&�ϡPc�4zbpQ�=���j./�q+�OǮ�����Y����7xiY��c0�b���ӹZro�&ո�T�ߣ[���DL�N�Aۘ��5�ZK]���tk��)-�����y}�is�Z��nKw������[Y�����ɻ�ϏH�_��z�U����#�%��i�k��V�
cV�N=?q�V����n�e��o�k����͂��7ջu�H"D��b�#E	����#��U�l���ݖA���^θa��+L���ܣ�yd�i}���`{4Sr�k�xB]8�l���JeF�KW����C6�֕	�.-�W�����7u�d^6	~��h�&��( R�}��K�P���榑��.�rM�z�Y����E��N�ș�?��~#Y���,�N�RP#�rFu��.]�=�\2O8KzFf��pKs���q.}.t�[��B"��e�o�~Z)L�{�A|�������}�n��0T�'Ap=q��cp�a����'�j�-���K��9j�6'�~6��ʞ�p{--6zC�Վ�����������hőT��{���0���6����FI��&�'�M��h�ѡ^fY�\H'|��b>cU^Y9c:d�����ݓ��~h�ډ�6�'E�w]\>�ǔ�<y�	�E���nz�BQ�~w2X�daՈBA W;M�a-��=�f�����Y�9��ÜqE���RG���@�z��g��X��g^���ף޲ԥ�*���XEܻ�-�G�����yU���U+Ѽ���Ӌ	����獸���u�n�
�A�*6��+~v�"K92�����M��{%<��ʤ>���Ėud�r*�s����M	��s��U��yr�;O�hf��V�CF��ZT�������]�z���JP�C ��c+�>� [��s��'��E�m�G�P�6��7ׄv�.r̈�pm-g�{�D�$����BTKK���Y@ӗ*�ةl'
��nI��6�f���� ���?7�k���ŸC`$r`w�����Pq��AN���'��MV�ci!�J��vd5.���7�@T����z�������NP�yX��f�,����2H?|@z�w �����0	���"z_�Nh�.��rw����+�bmM�����.��ܠ��x�ŭ�F1dI�nlސr�o}pLu�յI��97
�R�J?$���Apb`w��F,����Z#i��7[6�.L�bYi�`�/��h7�ވ:#�ךYD)%\��+�ƍ�Qs�[�`j�p��+�!u(�<~^U��1oc0̗��À��b[YP�3�x(��=C�jl8sՈ;4��� ꧙�!��X�D|��C�w֖hm�V�x��yF�א�UG��+�e����H�5���X��XZ~+�_�L��)L��W�&C��bKK���(ztHx��++~,����d�g�c3
���r���j
�	�_(�p�;%���M��9d� ��6x"h���?������T�R�%/U}���	w-[�9ܬX����}�>�&kO�����qf�wo��B��vfN�E�&k�%��Vf�� i8s��$&�^1�Rl���N-"~\��I���9����YF0�wL��S7�l�̦#�R[
z��焭����{N:�9��
�)3�ʴAa>�RW:Z����=�&o]@�
ˡ5w�2{�J����5	�ץz��Ld�u�Y����?�?g^�H�J�2��4�"�j�I�]R�ǰc�P�nZg{^̝>I�, �$;(�~s~���ޥ�޺�C����Q��
�n>��uB��&�C��R�4F�ME�>��pT�����ˇ���֏n{��N,K����yi�*/�pR�#��Y��+NeOS���ǌO��D������� �zb|�3��߅�^�T0[��O:���ӑ���,�Z$r�v��F1)�%9ːYb�᳌࠰vHPL>Z2������Zx����Hូ9� 5���[�}��(Vw!iT@��ӣA�>�q�Lb7�d\.�j�l�l]�� t��m�X�c/foI���S��G���]�͊�Mo� :ۖH&\t����c��F��s����Lݓ+Vv���w���`����#=cL4�bL��t����G2��� �:Ju��I����~��`�j�m����3�W�iRRn)y��'���̚v�l�=ʞȃ���q�<�m�3<^�=n �w|����:h¿NiI:7�x���*�}A�e��po]�e�R�z�R1�Aܖ8��	�q--]1��F[<��I����q����ڪ+!��Q(�Kh�'�A�9ͣ��_���"�L+��@��ڧ�7��Y=�]���+�����¨������
�!�Q�� �J@�}���L����P��QN���s�}m�*�%j�)�ν��]�k>���H��T#�;���v��� i|�-�!c��U[:߉���>�5��/C�<O�����=ϩv��!Z�Ǵ�0iXpQBU�W�'x����=�ߢ�E��b�7o���3ԍ���!�	�$�˜�<~")_DώA�e�=/���Y-�L�P�\a~�N�)͒Nd�?����ռ���1>����S��P����]>�2[H��c�?��p��*R�+��Ej^��q�M��8K(���E�א�-��6�����o���r����\��Y�%��"@�6�����=b ;��,Dpo�(��{.�]�H����������i�0����Z�};�n��c���n,8Y��n�3�x�g!�$�>`l�KY��	�JO#3�<o q�6��Ob]��)�<K�Ũ��U]�R�T��������ط�G�}v�"��8�!�J"&�3ɺ�
��b�i/��l�A.��f���zN��l�P<�6�M^�F ?�0�TF*���h|��"ؒX��kY����W`,,.�jlQ*&�&
�����wF�K[��>V�	1Y�������9���]��i���Lt�qI����na�Ť#�h�*_�A�W^x(��B�b�7��Ϟ�*!q�<B��і�"�Ckh�8��^��a1�>�(��VqA 6��p��-��|��Z�m��	?)�����j
�a��%*�&� ��;�B�
��H�d
� 0L�P�����s���4T�'���?��Q�0����rZ���!$�O����G���:�pk��[������w��J�O�O�㐿;�{��= v�S
�s��Zؕ�i���z�?�t?G�(67��3�.��
�:������ZCu�[,ۜk~�A~����u��.2#ݺ�l�N����R�6�I?5���ݭ�8y�/RlM�+s�tg�>�Q-�:��m����k�70���_حݫ��
�G���K�W��~�Z�Qga���!GJl�2 m*D)P�ʩ�L�z�=�}�����9I���􎂟6���V���d�M�SL�Q���DR��pz~_��B�\L�0A�!�ղ,}�=��-=�]|�y3��b�_"�}3mx�XB6���Jg�Pj�Ux8+m^�\W�{��:���|��R�3�W�uS��|9��\�U�¼��ұ�qY�]S��vQF�#�&w�-:H!�}o�.���4ʆ8��Z+܎�UX�D`�¡��:��{��-�sZ�9U�mz���(Ѻ��5 (���l@��S��XC��I311���ro�[�w��N����Vĝ�|秷��T"Y?,cx�� \��}(L����C¿gVegY�س�v��<�8��W�f��	��_���2�s�GDP�o>��&{Ej?����!go�c<MhB\���!�5z�4dWZr�wt.���ŗV�^�ZQ�'Q��I��s� t&Bx��ë ���%�/ߋ��Rn��a���Y��M��[�p�0����qf�Y����Z�]�m@�v�lHm�KU�t� ZM��U^j�(��,H3|1y3(Q��
������w�F�q�B��'��Q=���=U@c&^���@���,2XGޛ�Z���w�as��>�����QWuQS���56�����f�[-סG�O��A��������jgsC�-e���W|<[:�`ݦ���	�\`�Ei��G���X_�F~�8�	`��V�.{>�����3��
��*�pt��P�U����_�[��D����)���N��ŚU���OΛ�.��L��n�$�R��{�T�	h�M^d�,�1�!��;GZ(h?m�������O}�/_O�m�q� �1A|�\�'���|�吵��%��(����<����X�Ө~��K���^�ձп/0j���y�1jZ�� �VYM��j20H�>{��@�q0}+ �JKŻ�&�-x����^1��8S؆;��5�Ԫ���OR08��mśK^SL���Q�\���������b�&I���p�釋�̓'6��M�B.?/
r ����3�J����d��O^+'�������z��9f�ۘ��M:F1�(	&y�&���V��Wj@C��5l��?�M��E!#�b��F�],1�Ƴ Y��.�|����+�b��Uo�����Bw��սF��~.��`���lnZ��M���x�qH���~�w������q��`촠���������n�����l@��3A�	�ʵw��P�D�V��؜����R��]�}?v0%\�j��o����]b���
x)!Sc�3"�����V�L���W�Cx��_WD��d�'�E���A�
C��kN+׹C)��vx��Vh���/���^���:��p�E^�8"���xzҗs�h=l���86��X+��4�FE��_�㘻��r�*r�;��D�I�ǐ�y�m� <p�pEp*�2��kWIx�Smu�k\`��Jb�j����3�F1!����<��nC�0����:OZ�ij��ߝiy� � �Ǆ)�P�0��ia��F���S��)c�-�4�1{q��A�� ����umn
j�aG�j�!K�)8����$�N�Ȍ���c(u��,Oq�r����h��G&�5|4d3���L�X��`H�W�L��^$K������F��R6���]C0���<;��	90 ��:����C�;m����/Ȕ��&����3����]����o�o:L�B=��}[l=����D�䇷�t˶���¥�$��1��/W�fT\]_�X?9���[���u���OvAJ�<�]ҫԍe���b@�rXΤ��g���\�/�Y���*��f��#`s�i>a��~�*2����V��l@ �x�/J+E�=�b�]?P�:��U��x������5+�TM�27,W柙�����ʬ� �X�؝�ۇ�C���T���F1�>�V��<Ħ��hVN�t(� �y&����f�(D���Jf\��)�]���)�I<�^��<�桺��Nzj�ɻ�%��gr>u����R��x�w�>D7RN1tY�tt��)��.B��_;�gK[ǺF����R�β�NƆ�7gwT�5��9K�g�W
N�r���"���_$'���գGjv�	��s�4���!`�"�q2ّ���e�t�d�k@^�����ck� ����AG#,>@�AI���E(������*Fy@aL"|�R8H���Uɱ�c�S�	�y}d)G��.. x�� �~e%�'K��_�؅�&`bǇ▲I��ө���H�q���e��%�&�
�i�c?��85���++�%���5j�]����h/�M�a��s���f8"��;����'��Đ @�_���iQg�3�~�5Q�hI��Br�6����kD�PQ�8.���̨���by~�J,-,b�(�-v�|{�v���rwZ�\,��X��b�K),���6ػ�](hE���8f&o���Y�N�k����ڍAӮA�4����o�Q�|v��gJCxM0ϳn���)� �,��8���(Y�� ב	����)>1�H���(?�[��\��Ӆ} 3�������%r �pV�tN��T�2z���h_���ݾ�IH�P"y�ZX= 3B���7ޏ�Y���$�������!�ւ:_'���{����W��j�[~�����p�7��z�/lO|��b!1V��2v��aE�EEi���W_W%��i�8�*�!�kd�=��ĺ}�|�=�]�|$�����Z��P�,,
���`	�]�[�7jV�"�9�����D����52�(�&X�3bf�d{.��¸)���nc��Z�:��t�6lZ���ƹv��XJ�󪢺���b��s=T�W%�)'�~������5Y�րn�j)сr�`6/��(��(��
���*;Z��=g��LLf�B��W�K��g [�G�ic*����U2�B��f�R��I�^��A��6J8?���r�ʵ^rQ	�oE��ڟ��/wN�1Z��;�.�~�>��^�{���Б�p��� c�Z��@�+'���`F���@��x=\�$�)��$f��.�T1���!��^�	������rL]Lawzވ�?x8�� 
툢�m����jt`�8�Ζ�t1Qw���XܙЊ!R��7��E'Cn��I�>�p�r�x>���Җz�/D��̳���M�v�-�e"-�����Q \$�1z��v�������}F���"�{��U��� l亖�[0���K3�*�%D�f��bLH�;� �����>����e!��q�JP���QG�*�ؕo�c5!^�� 8������3�����z�R��Q��*�3n�o�UFr�r{< Vح� w��Q������$�\�$�=
]�_p|���rfԪ�3n�wO����Gg[�"b+/��I�������p�������`��h��E!��!HP��q%�፸���1ި��O+�Iߝ �}��oC��	�����'q�,����w ��z�6�U\C���_�\`hJdPP�<Z���"�X�:k���<૜`-�|�'A)MxN&�}L2�uEç�)����w���Wi<k,/��>�T�9�^' ρ���c�iȑ��pИ��r��9ӫEj���Uf���j}�n�j��&�F�O��C}�1g���-f���)� �~�u�x�Zj�%M� �h���������J��w�2�ڶ&%�ห%��[#ʐ�Y>���{H�-�)����؏E�0x�؄8VS�5�_E���:��r��T 6�Nh�Mb�Ǒhr�k����qBO�x��Ћ٨��įz���h�T�����i��.e���P�t���f2�B}�D��+5hk��j{�� ���e�x�[�������@�Z�W�>�:���NY[��h���˟�=�y������ߒ��<�{�RFR7�j���H�ͬ�"�Ǖ��/���x٭�!��$�TqC{�|�G�S�)Z��ߞ�S�+ݾw����ƙS�Ë��E�:+��>�&/��l��t3�@[EU۝v�M��(II��^�JC��o&d%u���ɻ��>r�Cl�N@����;qwa����W�
TdY�E^���z�����V�#v����Q|3�juJjfa�[rQ�4�ĹI0��f,=S*ǚO8�<Ep;�����I7��iX'N����y@i�\C��{�T��X*қ ��)����E��a˞�t�tjX���̷���D~��lق%�� �-�wE�Ͻ�3Iq�-ݳ��Gmv�t��iwͬ1�����A��W+�� 6(�N�~��8�q.���d�۫��y�j$z�3	O-��i�=�~]�Ը�U�%e� )�{�J�� %��h�@gKKK��m��Cs��Ga��A�������T�+V�O�����W�I�����A_�|p�Tu�V7��؏�G0ٹ���
�0��>���|^{����XzzS;I�� h�yY�y�N�\�.�1�<l����S%��q�ÄC����vİ��P��b!tu3c����<�Q�ȗ�C��Q��z��IG��%G�+
Zz�����](�i��er�������0�ܶ<�Wl�.���`뼳Ԍt���&6!k&vs8�C�C����~�S�q]�Y��Hʌ�%vRc*�}P�8�d�����A��SE!��������.k:��9�>͋�����������C�B�ѵD��-�R	X���7�m�?�O����W�xZ$N����g���R/b]Qէ�"�)�g���r;ۼ�Ip�;�4a/���?)G�t�Ũ�V��(�?BPF�O	V���T�J�Դ�<�6C��g����r� m��f����6����K���	�������fK����f 5X���Z�����O��uC\�7�Ry�K	�4Jڨi�3�߳���Eh���^I��i���)tP��u��qn��M�/������:�yH�/�o���/F�u�a
��T{�g�Wd�L�m�4���Κ꬀S�a!��z³(��"��bk��I�s$-��fYX� �WJ�]��ܢq�MXP#�t���b]=����,�[�BӶ�V����1�	���LcB���6b�hI^U�o���m���r�X��Y�v��'v�)%��Ag?"��p�e>��9��h�a)��(�8ϬN���Yѕ^h�z���{ ��V��� 	J�'m��-6��7�KH��@!L����C�P�C�k�3�"�rY��Y,ځ�*�G������`]�F8_x��a�4�ߩ�_��~���"��	���%3ǽQ�ಪĽ���T3a�l�Y�]�;IͮH;k28.�����\o|�l����r�c���x�P�������u����zs��f�g+p�Y���I>���tu�o7�ߏ�v��6�c@��xΏ��4� ���5?޶�A�8�LG��z����/�|!.��%æzx=o�aKqЊR��S[p��Q�n��N�P�5>C�[^��>b �I�^	���;��oo 3 ���uB�$�c��̇�ݢ���SXq��3c\$��)Pq���!�5 �c�ň�����[��݋��w
f���S�������^'�����"S ��7Vս��}�T�Y��=p�!(���!���=�tr���H�X�M���!F<ZrV^zL�(�1�!(͈	z��.[���ae�Ưg4)7�����u [r��bdb%�I����7"���vJэ��U}_�Q�!�����5�XQ4)�D�Od趃	HM��	� ��ݝ島E�7�#��j
�P�E��9a�V�W
�'��
|T���$-[t�������ǿJ�n^�թ�ȩ�4S���̖R�#�i-�~�^	U+�Z�,E�ڿ�[obJ7��93����D8+��r��%73NXP�n�?kd�6��<zlWI�!�[A1�I1�\�Ńb��J����}֞�H�p��	�
921x�{����DN�Yi�R@T��3v���LA*���rQd�T������p�7�$,gs�Q?��yO�&���ю�'G��u��z��]��8�R�
Dl�ҕ�?Y��z�2�d
�<R���4$>�5(e��0�%�2�5���C����g�A��8�[���!��
�8�cV{����qY}��N×�D�a��<"�/�9�L��l5���Ҥ,����~؅��0�m���4s������W?W��}��w����ųϿ=�y:w5x��Ott���+-����~|���C����#'R�%��ѣ`�+:�j~V"0����:�m�/�=~
Ͷ4�|�7z��@��~5Ww#&Ɨn7$&�"�%�-��J�q� ,�yp`�5���Mj���57�?z4n*���b�@s��4!Ȯ�V�j�J�r�㪴 �;U���>ׇ��	]���suv*�F�L%�h�\8Z����se��q�)b
7K�f��_��;�{u�}c����wPA�s��)��t�m�x�����'�+?�.��]!B��YV��.G�����FMQ�te"$Ϲ��[$�2�e?����[�n�4��<�/�IYR��f��7���xi����B!����l�
]�N�'�'xY|6^F���[��*<��CbĹ2�}��X�/%���v5��k-��k_\� :�P�˔�(J>M��B,�q1Z�{ɓ�gJ^�g.
�D��%��0��N�>F�/6������� �5�F�2U���6Ǟ�~���Q��7�_�sr�Οc�R}m���������r�ʜ�e���F�.���A��I��Hɰ�W�x]�zM_��U�>F`���L����݇�(=��rz�۞Uz����f��1M[3�S�.����f��d��t�K�u��߰�Eصq�#
�E�n�����؜�d���kzM��6g���*�|p�_�-ͨ���k�-�\e
��ìv�֕��̧�r�<^ ���O��;�tys�p4���Jkֱ�j`��'v ��;v�;0�o8r3��b�}�<e+�?	�]O`L/v�ONN����3h~���aa�	·�f?{;���'�u�W���劎�hqŕ�a�7����1@������I��W��f����ؤ.�Q,{�*��c���'��PM�o�`�C����+�!�t��K�V�_��*�i<r�W�rP��7�
1����:�Ң�n��Ȼ �{��[Toǎ�J�t]gH�������U���l2��K�� �V�s~��M�@��*�|�Aه��"�� �j�� ��ϊIzW�ƻ\�E�I4�0صޢ���R�˕So��y���$�D$Ze�ɷ*FR�~����Hp�nRL�3c�ⳅD2�ys�w�HX�^�T.��bok2����V"3�W��!�N}�i��>���]�)Z;�Ҡ�օ��.��̜b��p�'i����/�m���ɴ�,����;����iu�m�I�A�ʓ�?߆�kM�v����j>�:h����F7�0M.;��>�I���7���6\��Ƚ�������?l��?�F;p+ǂ#�$�W��rP���Z;|���$)�����Tm���;�BĿ'���Z'��n�N�_/�!3%�|��-~Q������y>0���|v�	�(U�E�y�G=���U�r%���S�'�Rc��Wwl�w'��*��Z`���\�Ӿ1�>e���
�����f���z�.���!�uߩ^ey�g���<����Ha�g<@s׵�۲�=q�Wo�+��=!jc��
��ҿx����7���vۢ���gO�����DDC�������8�~X�1����]��n��CT���{�;�}	���~^_�!	x"��B����.P�ԧR�%����qr�Q̺�.�r�� �R;�����.5�c�NER\���4&Rd����V�i�:����8��2�OY�o�!�u�!���s��W�k�7b�u��5l���/���H{��R�>�'���lgG�[VT%�n���hzW�̌1��*bs���ԁ�`4?��g^=�8�س�|�c�P����'�~�����j��>D����e�	�0[3.�q܁B�~�O1��/����4����"�}�
�#��b�f5н�S�a%���.��b2��p�{�R�	� I5�QS�t�Ox]~k%j����yn~1�AN����������_���)�9\�̚�X�$N��l����h��X����4I樌���3&���$��68���_.DE`Ik���c��W-�q���H���&N����S�])]��`a���#����&�u%P�0�:�E[���x�.��[:k:s��D���n���������4ж���(��#5Xz�E^�X��������=8�m &�4�w��Z�3Mso �[����7Pu��2lu}�*we�\z�	֥sZ��؂��p'��p�@K��1�ݴ�i2�z7�j�UG�z�v�Rq�|���ѡ^"�AրG�HM����r+��[�WiV�����}���Ԥ�� �X�t��FS l���ʹ����ol����z�A�.I`)0P���Kb.��+�dD�W�`�p���J�=|�֧Ac&V�9FJ�P�$x}%
�"?�Nj*�s��ӫp�MGD}�\����)�/�2����s�P�qpMP��f'b
d�弫F.t6�l��#eЫ�s6ByW���/��D�B0��^H�ʖb��ɑ��y�QĜ��с�$���������0����!a�G�.b��l#�w.yo����\9I/��q��+MrA�5�G�|U޻�F�q`�9n�M�2�Q��~���@��W�J�`~_��G��B�/��u��m�"���~��K���ӕ8t0�׷� M�*��*�^b�D�+h
��%��WM��WQ�:�J�Ƌ�c��]��U��_���=���ȓ&`�8P���cu�m�!�H�R0�ȷۉ�A�Z9VDKO��,5��ג`0	΀������x�Y�m��ڢ(��,{9�ٖ0l�_�~���K&ȋ��7R��Q�=D3j�E��N�R��]�[���J`�r�R$4+=H����w�h?M=���W<�¨�\\H�����:H 7:�4lK�Pa1����a2݋�Tظ_�zKޭ}���K}�5��_�6p#WKc�.*~��<~��㗟N,���ݳN�Sڏw�������v�g�e�������¯����z������P�|��'	�:���'胎�Q+����Z&"��Rl���1�z`/N�E&_�8��	.a���F�[}4{nZ+�q0y&���w���RȨ��%�K�}���|%��Y6��1��:hh��<�eX�m�=<00t7HwH��twʀ�Hww �ݍ -C�JIwJ7����~�w�s�s�Zk�3Ҭ�	^E�?ӂ�LLy[X#n)��b�oL�9ΣѺ�P����S�$M�f'���x��F�wu�+���m7�f��Υ����H!e���Y��i����Q�/Q	�]察�G�Ϊ��䕵R�PW�WHƧ��a[ ���V��fܗ������}�-�~����S����'�ּ����n������+���aK0��\��턁'Nb�lS���m��������82��qB!O�ˠXNl��<0kcy��Jq=��0�2_j,CE�s)����VIP���k7�:�m��#�_8��:��7R��:R���v?.Yo�]�%A�)�ZA�sӒ k��X��V���-q,�B�XCe��� �~O�0Z�ۤ��!|�5#}෎ě���4�TI3�h�4��>GT0��s�6z'D���}C��K��U
�(����E���ym�7B~���g,��g�N�иa�T&���:V["<|<l�|�Ҫ���^����-n4�?�9T��oZ��m^(�v"{�/;��~Jx�]S�~�����m.ͱ�;�"l�&��f[㲊!I�iK���!�������H��A��~z`�Ā�^Gi��`|c�w�0�{�(�3a�ڝ�Ԝr�p�D��r`w��XكR�X��[7
Q`F�t�e`*-k���<�SdeU��;�E��a�ɸy{ť�E���t���F�z�qnbc^>"e�=��[�Q�WV���<�W���Q��D������+��Q�}��fF��ze�)DG�J��rT�V
�gt��i��;%?�z��y��� uY�߼��S����?]k�8[��ImN�������>?�2�rtݚ��8����[9��V/OcJH3q<�)��z�Ѵl̺�=�,	l(x����I�����ˡ�C��	�y	.�����uiw��r@����{3��9��֕����g���.Yv7<7�*�֎WooVN�.�/�ST��l�-�y��iil���{�ì����E���@�y�ϰ�޲
��@�	'5��t8�����*�%�!��I��B2���'���~+�����7q�y��n�΄)iw/|���N��/���TE���|��h��-9"7�q5-5��'E��\+{��`q��H��͂A�735%�O`N�8����������t��p.g�/��6N/0o�-GS����V:��z��,{�5b�o�6A�%1M�0�2��[ݵ��Й�=��g*,�	Ë�Mص
�(9_ܷ�2՜̪:I���]�����H��z�o�~���p*��'B��%�O;X˃���v�WfßG���)WV�N�g�<���+/�#��c'-h�C�r/�C�7H�k7���>?���M�?8V��_*vd�<ך/��|*�د�X�G��%�^�x�ׯ_swK�c��ܜ���<�}ؚ�~v�<Ѫ�(D��	Η�ǩ���Y��@�lә��mʋ���0 �5@w��;C�fs\�0��,H�!������]ޭ��w��"��3O�Mh�r�Ƌ��4��0� �N��̥:��dI�~Q��7O{���L��ݺ�tϥ*N�� �[�<QJh��X�(��[�X;טA�<���b��ݍ0�V����У�9a~���.���9s�������+<V�Z�@�"v j���E�5�R�*`͒��!E�º�J��D��'ق�ajy���Q�M���@md�g\$)���v^���'�ï'fhx���밪����V����v�CY��ر�ޠCs��ѵH O�qڷej]�ݸ9�#�v<��h�����k����Ir�<�B�� Kǝk!gכ����˚J��ȇ5~'�?B�8�Xf��<T�#�f��.�w�-��{�(��~�}�:�n�C]�-���66H�'����VJ2�I���s��L�̧j�J���iw�$&��r޹쨉75��qX�z���𝦸4���5	���e�4�|&���>��vCb9k߉�ͱa��]�h�)��qJ�4�꡿yb��}#�TԳ�,�z�S�\��S�X�֭���]_F�8J�gOiU�.->�l�_��p	GP�9:�]��k�{A��w)����Y�!Z��J\~0�}I��ə���^W�B����Y�:�ӛ�x�[��*F�A�7p ��t�l�]b!�1�l>��k޻9/��P�O����O�fڕ߮C�,���oWo����([��\(��I	���:�|�wR{�����S��|Y���M�fa��iX�$]��eH��A���p����+���t;��K�S��|%�f��qu���N�dµ��!��di�Qvʓ�������ǌ�K%߅��aCvy�v�������H<�.^��=�o��%i��{ቚ�1bncؼP+��#������̺��o�C�W~�֝ԏ��	�x��1�c?I�#XmB��������c$z����vށ"؂�i~��:��,�sm�1��@[����u��2a�V�~�&���`�yD_|�U�[lYx���oBd~GH\�B�����j;�5���;��SY��*�d�'�h0Y���d�/�BC��S�����0�$3��f�_�T#���U����#�	�0�z���Үp�D������K��H,p��Qq�"θo9����D���lq�lD��7�"���3�w�&��Z������w�U�6�p;FY�>�9o[�|y��ilz�[�5S�㹎R�#_y-�и��:S��BjZ���;�0pi��^'\����v���b���%g%�I��}W��4�c�+�ؓ��D�RKH0P�	�k�l��$>�a�be2g�R�s�߷�q����ꉣ����?j�������!�5Yv�ca�@^�����O#N�����0tͧW��&�q4��L-/���|+�R�ͪ�i�H�9;O�?[m�c;Qi9�su�������LN�B�{�u�W��k=	7a ����3�h����{��n�����l�粳܅w����m�̦��Y��Qhcv��
��4ھ�h�z��~�aw�ӿ�}z#�8|K��J;co�w�w4'9p}r�S�V%������Gt�a�MTyHJ/vPhK/����'%K�Z��ʮ�N�+���xw�W8_t�C+�Պbt[��
�R�6����i���L� ^=����F~"5���E_��i�m?�-� �@[^�b*9� �$�����N�z"v�u
`����pFJd��&�6�C��������.����bT!���3`�|,�Yݹ����/]'�7+�/���/h�.���K'�7�[ׁV��j�o���\{��5B�ZAO�=Ơ��g��m�桢��'ʥW"a��y���uz����y�]�5���ai�4��۱~�����C��]�JՕ�64=b�g�j~��h���фo}b<-_��:�Ok^��-�}���V�ܣ�y�d��y����Q{��0��2�@h�����d?��w���,X湧܍��>?!?R�@i7#�(���J�'׮��zc�I]�\��n��C���t�&�E��U6��4�m�?�x��,x�ǌ*0>��\G��)�"[	w�b��Te�5W�����3�GP7�*�o��g�Ӆ����W���G"�7�*T�Y��&�NU��o���C��wmB%�hs�#�rC�HG�zl�T��p�
Z�Y���4-�ҥ���%�zz"N����)�Dr-���9\$�1�)���B��$�\��u��L���1$�n�f����)C�9��{v/?�:���w�=�mVb�S�%q�/Z�oZk'?���p����q�A�y�I̓����7P�9��o����Ë�
���O�Օ���ӕ�f��$����/GT�Z+�O��?�:�^;t�.y����9\�7<ˇ���hr��@������󭮻�*�f9)M���q
.����9�$��[��6�2�])H׀����0�8Ɠ����	҇vPe|w�(B/ n�.0=r�`"�>_�Er��I�
(E���2HFJ�4�%�
T�K4[���vo�w���*I�����Hg��>H60����Ϥ�Y���xz]f?5V��>�(i��|RDc��^@fRfS-���Jf�C��l$"3>�D�&�+��U?������R�?�M���I�̨K�ς��]ͣ��akmX��=v�{]�ׯ-E���A�^[B�~q�6��0t��O�8E��/;�w���B��Ϣ�k{+[ݻ�K��o�(OV��\�r�y���O����w��;�On�^���DQ�{<�>�ͬ9��^<������=����=w_sk�_:!���{:��kɡ�O�{��$���i�}g�����ɶ����kJ?~%_��^<�s(Z��߲5v���d1V�q�*'�/�v�'S�]:�6�?CbP�L�zlW�}�����G�����	������Y&6:���y�.�O��>Y�kx�0�Q:Y����bU7y{�<y�y%���-7�9rd�k��f��)9���j�x��rKV�j���jj��o52�|��ߚ�EJ��vq������\=L�Xh�����D��qµ�N�C���|R:/+`c$�"X�A�+ӂ��y8=NBP�5jV#�D�{ff+j
��5��ǁG�y
�� ��3+�HXԉ���6��X�������oyk��(6@y@X�O����`�YD�N��ќ�7}�:�;/2�!i%�נ�m6�b@)ɒ�m���_�ïԬ���J�.���X��������Y���[��Χ�� �i�	RY�i��F�I�%��c��ؾ��蓭CϬ�a^k���0O��aK�K�{dܸn-p�+����8x�i�c���n���q�(��3���S�d��%)ou%g��ӳ������?�}��!�P��i��!�}��X?43�6��I�wփv�h[�vtc��r_W@�Ԕ䬯R"�G�j�9��[����=��&�`�o_׏���[�oX@0w7PU�U��a�����4!�0I&jlk��(K��Uq��n��֓e�ۈf�2\9�&�U��V]#�XJ1Q=�0b:� Z���yw$��0��eW��&t.Y�h;���Mot��`}T�1�DxO��A�����u'E���� ���e�ke*pk��b.i쐩^սUb&m�`�
A�����x��X��u����2��[�m���I	fu ����%l�W}`�6r��Τ�\bM�0��B�6!��cұ�[.��:6佁��ި�tO�:E�(N�e��"W�aH�墤�*�:^����$���m>�0�0���!o�Ŗ�9�����"�3���Rڲ>���7�3Ұ�uO�򖰏�0�ֿqzC���W�
��gW�3�}f�g��_����s1Lq����*�2y���������������[4/.E���I�V\���az�}F���¾:7F��Ԑ�ce������V����_ⅿp��"%�֨=�0ޘ�ɀ��$�oV}��M =2��C .9�{x=x4�pb��o͉��]����A��L4�L8�	�.�m������g~f}�,��8I��,a	�(0R;��Z4 ��2��d���/���$��ZX� �
�ҵ��A�S3V0�+|����O�Q�a��dO�,Έt�ڢ���q��g� ����B��WH�������o@p��25�wf���ы.���!^`��Y��V��&�����+����s�֢J}�ɍh.�a�;"��t�� �����
K��z=q+�1>�.�5�G��{$Y>�<�F��ѕ���ͤ��*�r�y��H嗲��V����ѧүm��ϫ�c�:���� <����y�����"�}:��E�D3�S߹�/����Z����Ӥ�V���3ѫ4�\#(՘Nro{��8��V7q�����P�
��p��p�L1ˤ
K	���
�TBE���#O1.���Q+J߿aHVEK��!%�ˉ�"ĐruJpt��A����)d���T��*��I3�h�g4��]RĀ1[���h�^��/wc���'P�����
�&��Uk&�$ao��HE�^����N�\�>n�ɽ)�՝��{w�Qu#���nْ��0��J����� x=E.饟.͋`�a�ƭ�H�h���F�l�p�9"[qE����"_����p쩃�!����>O���~�e�_��,�Υ�r���3�UK�.|s��������BBW�H�����Ǝ���|���Ĵ��_� k�����&�V>���_�[��l�n���ࣦ���u����(	��Zc����ٱ�ټ&P�Ԅ�IʝY�j�+�yr����Z�@񿚔�#$����E�	�.S&�8A�K���;ݑcHE�������t�.\�[G��H���1�%��{�>�	$d~���ǡ[9����������3'��]G�M�L]E�]���4c���Y1�E���hP^��L����v1"��JQ"ۣ�^�p��s���(-@چ�덵M>�8=�XQ\��^�Qd&���,A1nY��$k�}S�?S�`��
��[㣍K��T�r�#Pdg�]E��&�@|� �N�a<K����*���_W��_�I���M��֍��Q��B͕Bg��g&�{帻���v�lstO +6F?�Н��~z�뛆kQ�,��]���ف��h�������R~eƌL������[���1Ob}H�"��c45���m�F�����-?��R���,����w��[�G�Kz�&�;<���}���	Nw���Nu�3� �9�9��q��3�$M޻�-����h��;4����o��o�+0�1��<�Ih>@��9v}ߛ�6Q���l׷B:��F��A�E��r��5�4��)�+����T���<ܶт��&Y!��)w]��x�Z�K?AJ��B�x��؁r�\�o�����{M8�Us���3`�!�G�E�������>j��j�y�!�݀���ё)\4򃵸�LԬ�E��C���l�eQU�-13D#�u5�˪B�FA��S蒤MQ�Mdt�<B�Z�4�G�^��M�{�v��D�zn�Db����m�%�A��?Lρ;.?ޤ���ad�ѳX��ƨM�|_�T�E[�x�9e7ʧ�78Z+�m���=�'�}��:^�1���Ĵ�k�37xRmE�hL��P�cxѪpx��S��z(5��7���V]!�Bp�@C��Z��Btނ|�f�)3"�j�1R���䯉�J ��2$�YDsn0���Ae,Qݯ�H�b��0�*ނ4c�&�*����A�q%q�r�H;ҟ#w=�0cL#@J���z��ɮ��!Hw����֛��t�G�j�����nR��ë��e�)�B�.q�ɝ�kW{�N;V�,��:�yWA�	���K�l&U�-J��{���2���;u��r3�����<a���#k��ۇ	j�.HQ������*_p����-t�0U�^�'�[p�]Q�=��Xz���O86�q^I=g:�;M?��������j��8���/��8r��c�S�1��tf8���4��x�P��5a���F��~T�
�L�'/�EM �Cm�أS�A��M�X��I^i��<�r�G�#��	�����H�NԱ�|Y��d��>�����W��2�?�O-�	�9sb\��O�t� ��`_�;.�2:�����y�܌�Ax<��z�w���|
��fsmg���q��Fz������0�	��RP���T�i��U5ӕ����0�������};6�w�^��I�ٰ���VVfR�4܍��t�`���+��Q��̔b�ߨ�'���d!BÀ�3ͫ�BͣT���MM'f��E1�ǚF��&U�z�e5oOI��Q�O������[jɻ�T!+�Ŧ�X2O)�WiG����S�7ɴ����[�}��#�ԁ��,o�g���ҍR
�$g�\||��~Ӓ�+i��yG�žz�� ��p�Wl��=���� (���B���k%Tx��P��Ʉ[��D�A��Ì&G�.�����>D���.�r/����*���"��!QŶ5�9�� ��~� 2h�/9^���hz'[��|�0��'���EO�[�{���3)4ȹ��?0����	&�u�Vռ�1�q��?�9�ּĺ��^7��F��|�X4E��l Q ��i�A��&j��6�5+�L{��� � %Cu�����׿_��[eY���q|P�U������(Mo/�
��(��:_�y�:�bp���&�h��9��e����r�瘝�h\čS������*�e��[~T�}�"骎EϝV�>\Ug1��%������E��Z��-��x2�oƻ��8��{�ԡ�.F�W��k?�	��a�a�8l��G����/�Y��y)w��2C�L/�z>@�D����߬q�M��q�?�Pڈ�Cy7����;�y��vNW��X�9�x���R�[�LG�8��A?�pB/���)���ɏ��&2���X�[��R�EX%`�H�𩒄k���[y`��c/.��5����u�3'?J_5F���^��U�os&���	ь󍨦E�m��=�w�(QK)$iHU�m\$TL2�neqg��V1��f2imS�u���5���X.]�f�pw��M�o�/j�Fp�H��W,J�r��C�K�gQQ-���M�R�7Teʊ�+���B�+I�O�+�)>d�5����߀t�,Nɮ��`|I8pW"�Wx+�ɘY��Q�q�W���V��(�5��%�䅷w�E���+m��n��Y(\�pq��T�h*�w=?Gό��0`Spp��A��zH��"U+�	p=QL�x�ߔAe>�`�2kO��q�WN��%åd�@
u���mS�o����Lg�����+�b���0������j���P� ���1DT@�?�#'\��8�I���Y��N�-�p}`�W�D�+UҘW��1���q<�"[ul3��G��S2���[U�^��T����DY�4%�� ��w��T��#|<�	_�*c�l�'K�dӱr�u0y6g�f�����\�a��
Q���89[�0�inI�#T�v������b\���s�o+������v�,N��I5� ��͢���d����9ӏ���"��)�i����O� ����#�9�2c�[�`{�=�j�������'A+�p<�p69�$����Cg�U8��G����I2�~�����7{�F���w�5S6�)�5��̾T��L�Ώ}|����h}��G�v��o��AS%E�V�]�;���7����@/@�l�!��[/8�R~w�2�I�_�!m /'3B�7�;x�>�������Q~���D+Gma�!zO�:PV��C���,1��ϡ�d��L����bxO&��a�
O���b�igI/���)����d5����=-zc�nh�������4��<�'���<4%	�.�YS7fU@������)M_is��3�k�4�M�t��2v}%$38��"-�Ga����&� z��E%w	��y�)��h �9��q�	��s(�A�x���������#��5M���{hs���q-ǲ���Pz�#H_�y���n���s�;qFp9֭�T@F����5m��q�1qer�*���O�^�J�@�8�V�}C2.�d6p~�P��� *uKꉏ�f��sXC(���$���������\�z�Ϸ�0�`C0km��B4����a(����dl�t�����R��L40�V��[/W�#�psjz�W�JVpU��3e҄f�ƹ� )�ه����s��q�;��9�c�l�VJ��;p��~��|W�9��ou����	��]gx���A�Z��j����[~�Au���&��CW�$�~e����/n�5��OO��5@o�'�1��0
����N��kE��2��@�-�W͠@4�x!Tp�O�&Z�0��u/�dE�c�������|�v�'�cT�-׉&p̏#R�� ��W�!��O$�����
e�����zӆ�#nc��X6�o��T��O��Qn�����^U`�Y�V{©g�0�W�nl�l�f�E{��Y���zN��U/�:���&Aw�\�|��,�J�"F���*��k�\��wJʷ��B��XMܔ>1����'2�7ˬ*�E����ID�}I.�ծVs���>�x$���F��g���
O�b���'�)L�,��\�!��CT8���^Q��9f������C40�x�(��������P�0'�}Q�-F�:bn�y6�����]x�Z�F.3�&A�[ȅ�B���<��k���fR�OV:	wd>B��  M-��BM�N��=��加b)Ξ ���H!͖����� �m�Jx�ku�hy}f�e���Ih���%j׎���_C]r���8W.Џ�2����_�m@v74uDU���-��نP�c�j��ʀ����O����"S!� ��P	b�1K�1�טw����a3B%3�$�+J����2�mعM� 	mk��g?:
�����*��C-M��[��
#��֧�=��b����4�ߧe��ʃ��P�cajlib��4��~N���vа��+$=B@���ws<�v���<M�Xn�Cp����P�!�>T79��� �X#. ^g���+z,����С��gҮ�0����8f��תN$���Fm)�q�&�f��W@��N�"�k��|�D0֚�(bM��f�2����1��;���U���D�����?��[�������@?�^�Ϳ-�"��	��;�
���S��g��CC��3Ƭ1��w�����L��i"�r7�B��5(�����g��`S�T揾���}R��1�2��_:�m_q(��m�U��)�/@�Q�xX��,���u[�pIQ+��?��Y{+l�ek'�q�e�����������A�y�H]�4VD�b�מ���N��"�7Rrp����`#�Y�֍���+�q\L.�)&���I֜�M}�2	�(��|h�:(�T�̬)�#o[��$�����_�p/%�=c|p�����tc�_Yj�qn���(߫�>��m�R� ��wX5��%�R�m�:DR��kϰ�@�6 �U��������B��^��B8X&
�D�-��m���E�= �㎭Ɂ��H�u��.F6B�
G�|��- >4(V�ES��u�zz�� ���lG �˻n�qCۿ��w`�&NA��?��b��H3�I@��t�ߏ7'+.�0�]0��O|8�
(�s=��L�a��}3H9fd�Mc�a�q��T8 �q�aR��_��: (��l\\�,�M6~�Ţ�%L��a�V)�B�I��H�P����G��\$�]���J*n��! ����@��Ə>5b�����'p�����`_���0¤B�&�V�_��*��Ш�R58�p5�ֵfY؈5�K?��b#\���S?��oH�T^[2Y�K[���6����N��/��o����K��L>|80e�=XEe���?#W��v c��"�hu�Q6X5��n͑�+O�
���p{��;����qVT��zb
���)M�9���Y���QxЁ{z�̸f-�#z�o+�EqLۺ���_<�t;ѺM�H��+h���ߦg�nn� �B�$|���U�8�p	����gա�{��7(M��w}ӌ<\˞�U�.r5�n̿ŅEw��UFCC��;�6��a$8��(��$���2��C��:.�v��rʬ&�Q%��nYB����)����3���}M�Z�3��͸���M\��qqSz��K�8�p����>~m:�`��w�vq�z-�=a*�����wֳ%�'s`RL&\R�N�C�_�|%�����lV��4@鲳��q�O� ���B�(�k��*�lݠ������"�?&a;2��[Ƕ�c�lRፉm�GɈ�;�0LS��D���"����R�ԝ, �d��'����HO3�æ��X�`O���9�",SW-b!��2w�h�y��q)&&nΉj�����n����a�4=�`ӫ��kl�H�!���8�����֨���Nq�|���=dG��>���;j����
�$E>����"�������v��rˍ�Z�'�2�_eO	�"{p虈r|o�2]!X����O3F��h/�z�`�;�ݭ�3�[��B����R��Mx��3��5qËѿ-�7��Y����2<�����lc0����|W`�Ze�4���M�W���K��|Ǥ�}||?s���w2��JW�`T��R[�?K7E%��6 ��e;��l(�3�͒5���l���r��r�w�t�tƴu�\ྜྷaM���@k�!�_�������H�F�w����(�����|��F���T����e�y'��۹�'V��܆���<�NH� D��8��6`�Zh��N��SXu iTa��+��C�����_9[���'\�]�s�
���i9m�0�K�Dq̓x�J�~�eR��P�(y�4��T2��3��!�WtWh/|$U���w��PY�� bn8.[?M�к8��1����&�[n��ߊ0̄���g��f��nd�g�iX/����<ýM������&\>�HD�"f��;<�i�k�W�hi}m�d����2*ŢtG6���e^��K�lkT!�#�|�g�1v���NKg�0�3ϋ���U�|f�YY"�N�(�y�{�����nW?����m?����Q:%2����"�ޜ��{E��z��^�7B��շ� *�g���Dņ���B�<q��يo�����~̈l?�c�2��2���ǟ����"�΅���0��ˍ}^m��ʼ�1�] ��������ArQ_8�0���D�Q�m(�Z#sk��	��o`��|��t.������s���w]?�Eۿ��$!pl�6T��?[�x��l��:֣�.���_�����?E��d��sط���m_�"pG}% L�Ąh�Ft�4�HA������`{�%��_�k�iF#ܚ��D2tp�^����L���
���f_5����#�[�"�;+���ғ�������%5�oK�SR5s����]z�E�8���3���������I�n�.�lo�k:�"�^[Iδ�H�z���o`rߎ�Nu��WW㿍W��·*���*C�!�X�p��`e��-��	^�<y"r<&%fHBetB�$��R��+�B1�E�����y��˧HH]n4�2ؗ3ZicuD�b6��4\���Q'�A'�'�*B�-�U��g��Y���h��CϮʏ=�p�X��{�_&"MO)*�; ��k�(����!"��[��6X�,��3͏�T=~7���LC�� x�R�����P��/ʯ�|H9���ֈA���}ϼAp�<��Y�ʕemPO?���ED>B�3POc��c�����"R~A�ӈ32��㏬(-�h����N����<j?Q�p\Bb�Gё%��m�L��_�w�$�'`u�&�'��ͤ���-���	��0Thm?A�*�*�"���po�0��*�W��$��%�#,�V*�M��;�Z��Կ&Oq��,eèǱ8.Λ)=2�gu7t�O�\K?�!�\�U��Jw��1ls�Vx^��	�d��Ðd��p�~1����B1��܀}օ+b�`� �'~�j�}�p�����>���l5eX˹���PBD�E�"�!��r�(��"ݶk�쐤T2��D�hI��x%t6n/�n��}x��+8[,�o���H�k��1���U�
����_�nrN����BP��|�>C���B�g����,�,'v�����r�uw����T��7��cSB=TU1 ��&y�z�P�E��b��?1j�̘�͖���a�Y���S�ʂ�y���;�A�J�����v���E��|6���
3Y`,����Y���1�_U}�	���8����B��9���{뉼Ծ��jyL������E�݂�b�nM*c��L�K)L���O�	yh!���ìy�`7A�h=t�k �(�i��M�?���^���<o���W��D��?��Wn����#ʀۂ������?"}�G��e�s.��OY�	6#ϓ��һ�dQ.Lxp�]5Wd_D��h���!��+��l���y��G�Zݹ�P��CeOW"�?�,f.�KC�w�XV\(�d��d�FL� ��������E�� �.��n��1O�/+=�\�*���P����>oȝM�x�,�ɱ����?ć����ѩ`ÁI�?kk�r()#8�|S�e���Hb��v�Y�Syvul �Y܍#T$�Yy�<��bHɜ�(�$�����CO��$�0��Ğc�qb�}0���/��`�"DaM�74����nc���1�����z��)�Y\o9B�O�A���N��%Eu��ҍ��T�<�{N�v�qE@<��}�~�5�������S�S��*G-J��KJ �u��l�?��8�Nf,Gx�Nr�F��v��N?�ޥ��K��룅1��jN�u�y�]� �{0��&._VXWD|�\�]�e�/[3E�>>��޶�]�%�6	� ��`��ҝ���h7��ҽHo̖�ɡ�*��R��D�F��%z�� ��� ?;	_����g?8#�tm�rN�Ynk����{#/f�~S�;��6{)�OJ�H�k֍�w�}�Ν��6M�a���xF�KI���د�4�95���E���1B�/Ncٿ֍�ڐR�|4�?ʩ��6Z��}�K<��ִ���h튑>�`!��V�*2����E���U�	��)S�R~�5�7��}?gޗAIK�?r���g��dЗ���z��j��l|a��i1���r+&�'�}/���վ�vԖ��>=#��<�C�	*��n`hخ݊皿��0Z���~�)�ګ%��q��#�?-� �X�J��^����I�i6W����X���e��G��q���8߭�|�3쒢�9�[�Ҝ1q=�6���o`$q)�W_�Sr�w]q��BrN��b�2h�8 m�:"��*�
�K�)0����I9,[��=�i�Lp���w�������&	��l]Ew];�[�`�`H�h �x���_Pڋ<F+Z Ia�����׌�b?�9��a�v>��37g���Yr_9T���6�e,�.�5��� A�?W�zViT�%v�2��R0squ'gk���b���!-�e��xk4uiE��3�$+ko�!ubGOΛ�Œ��ae�j�GӀ����eb��@Hw� ��2��d�i��1!���\��aˤȷ��1��#�,5;zz�o����V}��j������T���@�Ё�9`�x�}p���H=���Cp��h@54����^�B����7(��2���ݿ�(�o�1���?�e[�o?��(�(��xج[[y������E���􋄻8p[���x�&@<(���(C8��#�Fm��P�L�0���O�oV�&��M}�I��7��}z%��}}�.ϑ�O�I7��!k��{<�D�e3�l�I���������6zz4��y����vK;��A\]��
����#9E�mQ+);�'V���]p�"�h�<��Z�1ʶF���B{V��/6�v�T�������6����zń������)MWs�
Oc���O�tNM��'�ݤ�dځ����<�\�����$�d�,:�K�k�q�|��O��딛��ż1C�=��&�L����&J�'����Q���u��W�[�%��j5�*��+���Α@��g�xG^�j	�R�#hid�Q [�>�C�?�r�.���g���>��mz�v\�bYǉSQpށ�O���z��=,8�G`���;a�㝭2�`H�S5LK!����?���	#���r�3L����h����.H�^X�M�LR����h���Ɣ
O(�S���K3��'��*��D\����&U�E��E��>����v.��]��Zt���I�-�Bh�@97�T�����$�[��!���N��>�>E6Yg1���JW�!J�J�G}B���''
��n�0��'��8�0�;�r�8�0�:�`u���A����aZ���-^��!���4ҷ��7���qUG�ZxB����ԯ�}�l��-p�)�zN ���l�W>E�xo���?s?6<�������e�X�f�~���%��DcT��r�KJN�ɯ���-���{�y��>��0�Q� �9��`��5̈�t�7�4���NT�'w� 9F�Ùʴ�����I=�A˲�}A^!!,�lK����Ik�E�8��������X��|��<��=�L�
u� ����}�"����Li�Nq��x<*���¼��+<�<���o�N%!��G�O��a�u�WRs���!Z�)�>��7�<e�y���*e�Ѡ�����r���!���z蔒n))iDi�R��c(E��	�i�����e�=��<���־��ӣ-D��)�qd�����^��'��'t��E�&nbx���i(�H��`��aU�}���)�M�������[�D/�ʵ���7:uif	n�+|�jt����!%�)Ww������n ��l�@��X<�uG�����n���������ܦ�*p�a~����LF����u&=;�rWS�&e�7v�t���yH/�8s� �
<�C����8��z�q.\c������l�8�b}6��`,� !���SY$�����`S4�?L�c����r��rPao�BY��߹�^�(��)���	�<����:Ҭ���A'� %���Ñ�b�eL&���������5H(� ��J��3�x����l�ƒ�@�`��L=gͼr��5mGq�n`����L�Q��i���OVL��Af1n/W�A��e,�\�Z%F���/��vI��[J�Vv��
?��?���넒�"-�F���{���mF$Y�
���`�+�$q�慝�[�D��u�I�ć�$��)0$i��]�&�·ݸt?��Ѵ"������Ru�l)�ӗ6}���ϰ�ι���#4���M�3��<s�3�]�aב�D�E��/�U�S�����I��f�[���h٫iuR'�YwҨήl������U�y^©��v��1��nC����8��j��oxT&��`3��D�E5c"K�޼^���"�I��-�����;��A�g-�;���jW�����4��f�J�&Jɶ�J)���+b��F�MC�����vI@��c��<K�a�QC F� �=J�(?�o\A��e�{�\m晍��i�kjT��%�c����zc���h"�Uq?�,�О�+AyD_ER���x�VCN~���t(�Gg1vf@N�:}���=(�=�$��I/��*,A���S�es�Կ*�I-�ɇ�i�a�⵳�2�c(Y�zY̑�J>v��0�hgu���W�A�����`z5WA��ӻ��5��#�y�5+��l\����w�	���s��ǲ�;o]�'kL��
���Ǆ�٬���z�b�h����y~~ˠs����l��������޽N�ǏeE	�WP���%���N���Imť+b�U�,4��^��Ԣܽ�_�鼅S�>S�l*u�ĥ��މ���e�}�9�|�˿�A�|u(��U[���%�1�wA�C��_5]2c"�3��~ID�EDL���gaQ�'���@�{WH�T�H`'nw�����r�]s���gݳެZd�Y��'>�I?�]S��ĵ��J�LѠ*�L~f��W�\-#(�ھ>�2A���-���jH�������F�Mg���p]ie��t���P��	�e?��;�Kꩴ,X�{�	���CzQ�޾?�O*~E-�U�ي��ɒ�i1ne$M)Vl��ĝ�\#^��\#<v��Y��_���a�`ק�[��u�Z{�,X�������at���Uc-�^�wO�g�����toW:1��^<��G�0���1PpV7FyҸHRn�T�=����|��ɛ2U�qa�kL|a]:�w⪿�9��T6���v�M��Fv��F���՝��s)N��8��y�H�����ܧ��n�����O��l�Q,u� ��赲��]UO�|ٻㄷ]��J�AR�ﯷ2���0G��s����.Kf�󫺋�����T�k�_�EL��?��Ӕ��}�x���ƽE�����W<2�3�C�WO�:�:�8$w��U�����w�t*����h�����^j;*L�.��RE�ك���znr�iNZP�@M����
���,S�bM�,"�{�9W`Ti���%�a+��_r��Սgq��\��k$&���\��c��	��\�I�Y '��ӗ=6kM��ڪ$��ANz��4��6������i������xT�] �q��Ȳ�>�܂��D�����GQ��Q�6cq,Y�*�{���i��*�nᥦ�z��ɍ�/Zq��ފXy>k�0�4n��l�Z�Iڈ���&뼓���**I�r@�ԙ.��C�����,�Y�k��h�#^��(�W]eOM��T��Hk��Y�
89DE���7��0�K�j�3�/};�A�����<��k$����g$?��t���@+V��[w\�@l�l�X<7Œ���a��:7��"���z���#��T2������c�whᯉ�(�EU�s�p�8'?+��!�1�_	b�^O�6���=�i�e]KES�^���%ݔ�tcq��%&��D����"�P�A�>������9�k
�!�rl��Z۷�A��=�B�����-�2qg�W�t��-�R,�t���#�R�+
�.��팇ەG����g��H-Ɣ�uݝ&�俯>
F�0|���ol&�IQ���{)>/ݪ^D�@��Ā2�x�O�^�߻�!}MU�o$��DB���4�J_�N�sK��,)�ț2n{ʹlI�֧V-�-/�N��!���Y�9��Qu�C�<Zm*���-ޙL�bu2' 0�{kz���m�Ʉ��{���Ԍ�\�xU���3�Ք���a�A�j[*K�v�I_��L7�
�
�b�t��t"�!74��oRW����/QQ���B ��e1�|�m9:��w����0�c%���<��nM|�-��{��w��Эt����%��#��Ubۯ��	������W�|���b0M�M�E[u�&�d1�.|A�5��>yK�J;�~�O\��2
�B����|׃���N�B��H.����ɠC������jo	�3$�ρ8M�q��ڶ'��o�̦�d�hȱ��.�+lb� ����~4��H���R�uIci�~���&���X	�v���&ϩ�*Y�~d��+�S1�rVS�� �#xZ�l���SH%��j�?%��e��'����w"o�Z�2���J^t��^7�c>�VS8�@T��N2�t�8�}H0`����������]�֩�gF �Y���ר\}�Ab u	~T�Aw�Pւ�������e?\�����[)1Cŧ���̓�k����g2#�^4��� 㼆m;�`�Q�c�M���R������^8�U�JIm�HkC��O���O?�X�R������R�,�q�Hix_.����^:Y��������b���ts����w���s�Nx�;�2�	vQ�#���,!����*w���kw����f@N}���7�����7��̮�K��̴DשҴfPan�f�á4�L��ڗU0�w�Mu��{��L�rf���.*Ze�fk����O�����͔�
�HS��=�M����	MiԊTt6��$��~aηTRGk�����0���85=�}�Ƿ��%�o� �Á|��:�ޑ����GZ���?Ŏ�&p�MCI����hW��<d�D��V����l�'��{��>���S$�@R+@}�񍅜����J(���K�j�S3򚡎���S��e�q�nUz*~+x69��j���l����K_`M��>���:�_s	8a���j9�I}N�kյ #e���_S��%�zE�Sձ�'~�ҹ^� R�X�(����3W�+���NIG9[N�S^�׋�8�f���re��V�*�"��篜/�$�;+VC���صr]��(���zmQ	^+<�E���fE#�f]�}�;���Ξy8F:ZЭv%)`��� QDl=���Q+��S@\1�o�|r��jL�**���-q�Bb�.�l�'̺�M�� ��Z���^>Q�Z�7׿�vqXO�ܐ�o��=������B��)�E���.�u��2�� ���a�X�W�x5OR��!XƊ�?��t'�NG���qm�U=������w����f�6���B����]�	��G��^��ǂ�e��/��L���(�VgN���M�<�X��lh���%�����9�b�=ʵXoi4�:*^cM#�(.���Q+��43�] ���ޞ�!y��(G�?���c�r5��Fh	��wɌUkS���w+T	C�����;��^+�i�a/�Q��JD�S",��M�)���	:�,�����s�N�(�0���Dp�,�Q��4I?%Z�?Uy�$�ڐEU�~��1�L� �mڱ4�� ��wyM7p��!-�1Q�[Ո��"u�V�P*q��q*����1���$����#�����Yv�m�"i����_��d����'w����_����P��!Q��A����2£���:(e7�;�eN�h?؁��Ԉ%v��р�$�{5:�=@O�P��w2S�t�{�3-3B(�Bc���y���5�3��J*Ƌ�q3��@\�`�s.
x11�ջ8�ő�����]�D���'v��r'��d�z�5����U���B#�$kء~��(����_��a=���o
��<��
`byԍS�E�B�W��rK�M��
T�mz������$��j��\˷c\j���9Oޜ��E�#�!	^Z�0S��r�a��;{��ah�K�ߎf	�w]o���z���
��Ia�~HWf���	h�$o���P�/��ǟ��r��j�[��g6����08K�F�243���<O����x��jS�􁪶�-�.�>z7�.�й�Q�:���@zU�/�Q��8n엔��qf���
����%�uu~R�x��$���&��_�A�U��� �U���c�{�F�Y�,.��̐��܁S:���r�]*$ܥm�\Vk�"�+7�8k`�F4���a5����I|�F�x &�,ǥu�?�<��K��U"�����F��W�	R�#rs##|���'�\g�{!(�K��S���\��麟�����˟�L��w�)~eS�8?�D������AfU:..��7�5@��>���(!m�
�(C�A�/�2{��!�GE�E[ß�(DN7��z@[]�?��Ƚ�A6}f�oO~�����K���'V�e�pg O��2!Ϋ+�X���k# Vˮ� �=J�,���̵F��l�xQ�x�����}�"��z��&-ǧs=Fw�I�/�����/on=���<���q�Ku�R�R�JHN�
>%}B"g��]ߟg��˓(�����ʹ<�q�K`硝Ѫ��Q%p�dvӢ����N���W��	|O�1��G�Q	�=�,{�M�/Ķ�"x@�qS�����x�T��+����ѓӪe-4,�y��c�.�6:Y�sMB$\�Z]���J���/0�B�3WbJ=h�:	�u�tn���[c�R?�aO�� 1�E�Wra����N{ӥR�
��UB�K�#|�3E2��TS:�0%wQGW-O�+Y�z�n}�1w����+�@���?�䖹��'�[P�[v������x���I5v*E���P2���nmL��ཡ���̀�`l'?*GG���(
=�F�9�}pF!�4�a�Ak\�\�G���{�Z�l��ع��9�lԫ����LR���".��su~��º�v&Ԃ���3Q�Ni����kƾD�YJ}&��t�S~�'�܆w�l{ƍh��1�qU7
�?S�+��ti�9ϲ�vx�N
>@2Vn�Z���s���t��:bz��7�-&\�ɢꬺ�����!	�@:=?h#N�wq�����6Wy�X	�|���;s���NIP�:���<�+�&���b.��m2'��݆��,`Q�*��N���;��	+�����`��^w���5J��9��xտ���ܚ�,K��]���hu�<a �8R'���x����y̶����?p��M�i;1��$v	���9�,�آ�%B���2�R[.�OH�_���u0����ھ��܎��:ίO6i�EI��쀚�b��1�F����D����	�˥���?�ܲW�Um~k���FϩD��'��9~|c�`��13T݁����Rz?�K�MWr���6��H���E��^b�x��U.8o�i���D���ϭi��Y��,�����{η�&��n�j^�*�7�pZ�z�`���5G�;7<��X�Ago�*�aؖ�����!r2��C�Tݫ6��%%i�$Tپϥ�iu"4�m���6܁�X�b�����O�j~�����bdMw��a���������G6�����⛾�>aET[�G$�on�8X�_�(��5}	�U��y%����V�s&#2{
f��ﾙ�,�Ҵ9S������ĥ�9:�V�ܻ�\�+0�fx���1F�=C(��4�x%="��x/��݂�5΢�Z���ќ�4�j���>�?E��W=
M){Ard��!&6��B�W΄VV`�NT�(�:5�����+>��잘�a��븋�Z��l0g�Ơc5����S�hl2V׭g�ݮ��x��+2�x�Z�#��j0�V�9ش�������o}�W�~�|�?Xl��z|�B*٪�oR��o (.*�Eͪ�띮�}����X�`Z�r��b/�3a9u���޸��#%D���b+;s��%T��~�W�d���4(�}���o5X���W��-���$[X�V�W.ے٩r_w�r�\�3���dPU��V��$��L#���,H��i�4b�F?c����b�������z���q|d-#�(�
Z<�o��p��X��o���l*Ԥ�@���P|���w���,���S£u�����HX�P,��Z�G<�1bŶ�^�{f?�������a�����dt;��}^���$g��Đ�|�hX����"S��w-��;q<V������ɥzp&M~h��q̷jsIv1�-W�m�q�87%X�uht*���11���(�k�Sq����`!z���$4��8�e^�%�����0���*�قv�Rwǽ��땠��v`�ٶ�cg��C��'�/�l�¢j��&��ǻ�����_o�h���͠�VV�%��ωn��Fz�P���b���L�eB+�$/`- �,��;�<_�5֡? k�^�{�m���O�Q�]d����^Q���;)obΫ�S�9#<�c�H��e�F�_J���h��ȓ��;�ߣ'���F:r
3Ե��}(�c�|�=��y����+�Ho�[�֑��(Õ�&dn��&-n�&d����\ܞ^� �[-*�d��TS�+o����#�e|>����)������t�M�y�f�t������x�ۋ�`��K�д)r�+B��e��lcF�:�.1Zzk���	��ɏt�a�nTC�J ��~�T�ި��GT�mS� Q+���*UɆ� d+h`�MɂQbtpؼ}}ڥ-e����P�-k�	�[eejhi-I�1�OƬ������Vh��;6qx�[����̠ၶ�E*��1����-P�,켅��r�T,^�U2B�j6s���AٷW{�k�+H�s��l�h��ڕF�M1���bK%�F�(1�b�e�(��䃈܊2e�#|T�UG�6��F��D����!D�?s�t0eq��2#k�2�k	F�SuLc`�U�!r��ֿ�4�;�wF@lN+�H+ѧ"m��z�`=�*}�6*�O������Op�Z�E�+�;u�4B��f��>��4�!5��
�
�^��$d"C����?�?�_♝�W�u�p�	�p����7��T!4�v"VK��Z./
�/��j\�;0��~Z3*��@��a7��[r0�`r	�
�:�����z�AUN+�s.3�R��.�^p��r��}:�?�V�
���B�<ܱ��)�$UXۜx�aU&����2�{Y�ZI����r��x����y���h��Bk�?➯\׃i܎ߓ��nHKDS�v��8�h|��vp��&�>Ɨ�2wu�A+?'��E1x��r��p��	I7��=��G�to��(�d�6Gh@h��g�O�PuVk�E�|� h�{�34�#U�g���*l�:��@%NYpTc=�N8Wc���ˤ���,T��pF��6$	���7ݐ�R��2*j�y�2�(��cR��(�$���0)@�������:�|���pn�����Q��"~���ʉ$FM巃��1��*6�a�����c�`��uMG��^�i�����*����:�w���>��5#Ԙ=�cg�Ppu|ף�s�H]�]�aO�d�'CR%�p�EYf�!Dr%� t�C�'�􉿅D�(cb�̐ x�nY1O7�u��קB��l�Ƀh���Y�3/-
p8�ս�����(ը�������"@�L1�6߯A�*�O��rg���� ��p����z͡��ņr���Kٕ_\�Ϩ?<1��_�����<ы���%PR.�B��ݘ��o>% ��'�����)V�`��@��P�)W����\|��J�����d5�z����$�g�h%����T����9A���C����\�{[S��{
�q
r6ĵk�c�������r�����C�ˀ~�ZAJ\�1@��Ȝ� ($�p��P�
� q!�FD�z�r0���'���H��>m�����f�џ��^�G��=)�%�kf�2�a���º�l����iG���k�!q]�,Ѓ4 ������$�G��d�Q�:ZD�V�4/�	e�>I�'S�r�rA�aԦ��QC��e�V�2W���]A]`��>�PNIV�k�^m!�.!��Zf�)�Z��=�^�<Z7@�#�& �a���� �[<@L�3ӵpPb&[���c* ��55�[{�]Q ������S�L�w� Z��mi���7"b"��4Dˡ�eѡ(�NG��L�M+{���T�y���G�A����)������n�\b/;Od5�"���z��>�8�{�Q���A���W���!�W�w�;�=�& 2:ܚh\�l�@��(kt�E��Vh�.�.4H�u��"�|��}ܬ��:�h���)Kd��<*P%v��j�淩�4��l�!dg`��]�b:�����y��7��"�n%[�m�h˼�����{�Xc��J� 
�d���20ѡ��$;%�PpAJ(���
*����s��r��8ni�B��X�cU�<�ꫭ!���K��vt+&�:�nl�Q�٭�?t��*�pF�����{��g��~�Υ�Dgq�a�X�n��
�N�aL��/�C5�z�l��/=K{\oD�cg�v������m�ګ|�v(g�	Nwf�� �D/��
8�M}�������P�iT���h.�~G�ѱ"ˇ8.Gʅ��n�~j.&S�p++�K�x4�Cb�A�@F���j�P�^���/�R����5�gkE	{���.K2��?]#7���51[&��r�bԥ.���:��i�q:���X"*�& �TǊ�L��T�ű.q��s����a�@��0��w��(�X�S�{:J�'��|�����=x)�l����%�����p�)4�α��2�;׷�@3��Q4�j����Fݸ=�R�S�BRd]�#��u���� �ɫ��a9��_�?��$�H�`dk4Q�l!�޵N�`u������f-���Э|v0ѭ��C��tn)�1ڻ����i��(��z��ش���;����5��H�dZ-��˂O(����(�h���ɸHG�R^�����o�?cMj�:M���l��1lI5���P#�Y�|�"��k�>����?TL(�C[�!�`�Im	0Q$`R)���ɥ
�F�4��Q�����i����:$M�;~K	с��T��%v�ٵ��T_�<�'T����Ͱ�dlp�O�e���R��TtP��O���IP(��
�a��1�!�Mρ��1*?�ͬZ�%W�AYO�v���f/ͦ����T,3@�˷��&r~t.t��C,Y�:�U��,���F�:%���mR�q��T;��@.4����xRtu�d�4���W����Z�|'��F�k>��*<Xn�ƍ3Z��O�3 �Nn�)�Ly�u�t���,s,s��VƩp�Z��R�.ꍹ�����s)xy�F�̋s�濥n_
|������hR�)�i�J��-��;�꣋�.N,1X�W(>w�9osW�SxU �V��?q&>ț�����h��LnO��E�, ��`Z�;� �h%Xtp (��V��B��i�cU�GU�d�����o�
�
��Uf��8~�6f����2�i<��x.�b*��!H _7�ԃp8�A���Oi��6��l�E�j�K�3Ϟ�ivy���^>�f39�Q���^Om2�	Hp�j�߱�U��Ο%�J?�ƯJ��)����E�rʶ� �T1USj��d��H��̰L�ۡ3nO��h���9��N}�� Gjqϟ���idX�Q��2�UsZʿ��f�4�� -s��=�zko�=l�<���x�@�oxC�\-�E���l�da������/���Ry"T���a��*�i�90Q���.���d�%�؈�c���|��u����=!uKL�$�����V
�����������|i��YNP0�������cT�^+
:�Ӕ+ M�
 �鉋{�m���$�n�C�	���j ~������T����XN�ԧ�O;F��'��Ĝɣ�ߚ*�d^�Car����r�;��R���A� �  �<�+]]�2H� p�Y]��������+�8`����C��������Aӎy{vJ�qn�2�\�|
w+���{������V����^ LY!�O%<^O��I^4����W�?^��ߍ��ܝ\����{31(��N�7hmrQ����:�.�ԫ�'镼r������:�n��J=�ĳt��t��^�*0�dV-�'.�p����֛�y����S�G��Ψ����͞����hEgcsu:��+�@t~�Fܭ���P%ÍQV�V�l� ��I�np�x�s�v��q�PW��ó��T8��%!ɛB\�'�qF�tz<�xUq�"��Î�0JQ3O�[0_߄�|1�h��D�Y�
�
 ��%
�����9{~�k���Q�8¦����F!c+���K&�[�²��,�ąa�ҽ`9�B����Ö����$Ÿ�}��X�E$g����_�#�'x�whxs�R*�HG 	��c���#M��Ky�LL�ͻ،yU\��nB�Mg����kn�b��%�f�x���So���?��nd�>.]o-6�[��������<�i�F$z�ӧ0q�L��1#�D�xދp�,@5Ҋ�ڜН+�=h���'$�x���\BR�m`Gb{]M�8>��8K�j ���C�4߭��Ε���A�y���/�n�b��BҜ1�U�0l�����H�Um���ںMI�.�$��S)�@w�8�A�W��j���������:�y��
�*��hWD����b�M	S�^*c� LL�ڲ��)\CG�h� 
�؈�C�f~���|��'�-�k������ޕ�j��'
�U܊��-;��A�]����k��]BZ��.�qp��z��RM"
ٖbd�S��I�A��%�-�eG�L�ț�H���`���J�B���s��܈��J%(ToلN^ �����������r�h4Z��ҝ �Ş��2ae5�+�;N�}3�nv3k=��2]�ey��+�DLc4�+J��{=��,#_�JYEefBJk�(�[�oI�Ζ��[4��}��>�?f-,�h�	&��%M͐�.��8U|.1IEv�"����{�:�{_��6�o��Υ�����'6�=z���tI�0��G@�yl�|(���p̗Lo4RxEE������`�M��|��"���3%V�=Y��O0�-P:�������-�Y���a��q��+~���ruśB���e��ǉU���2,��]����'O�����\�P\�Z�S�Q�G{e����ޓ��7��|zh�4 �tѕ�����n�:����G���	27)l��T�N�[9ƫ���%W����y)*p�ݷ:ʣw�%��_��&����G��\�Z9�qq��r��c�~ZJۼ���z,�5 �s�$hBQ��T���"E�O�Q��qfa�`t��BO�Y>@��ٺLN��0߽6��a|�ľE2+X4���#�;�xT�y):!=	���N��}�=3mo�c���@�ʗ��p}wy^f��,�P��<M����\5�[�o�������-��X3l�~D��GiM��O�i� �=��Nq�	�y�8���|Y֎K�ԇ�9Ó<vW�_�_��le���s�]fN�
k%��%9����)�Uy�谈�2eo��K�_;�	5��1|�)ΐ,�~����g�����	�@nM:�P���|_ƄI<S��:t����� �LQ�[�r�����(�A$a������2�d�a���
����s�����F�hH�Ոu5��%1j���I�[��gX�He����g�ڻ��Y�V[a��ZS�9jPg����)��-�r҆���c���ĭ(>c�oL���Qk���x�4^npק/A��e�6��,X&U-¼_&S�r�������8ؓHk��/1_j����%K���+(Dh��b|�C��A��G�m����Q?��7�/le(Δ�]𪷓~ܛr��UZ2�(Z�hW�q2��Y03���a.�K[���%��ڗt5���Z�z��@���g�9]K]��.)�����b�eSU?�J���t��.vSDa��^T���C�ϰ�\
'я��WAq�&f��VJ!��]�T9tBf	���S�Jg^G?� ��g;����=�.[�3 ���B��=�w�Tu�/m0>㤿z�1�\�%ح���޵�v>5�=f���	�d�L�4Qb�U��*jw�-��0�����#"�{6&�w.�� �#Xm�����p�O��0�#���g�N�"j�+c�^��m.[��BQ~�p����������j�ϱTlV1*8�D�ZJ�,<m���Kӎ��`�,
؋t;�� ��"���@rK�7���
��+)���G�����T��Q�jmKh쓧Sӻ�&�-}|f���-��B���xN������>�`:��5���mf�Q&gJ�0���o�wc���ϧ����̄���**_��E�XJ\jX�'v{��r��ng�b���(��n���=Mt���	���vzu�՞�_�*�ί�O;k��Օ9C�O.N@UN��E��rD�[���~��J`Q�Un�$�f��m7l�6~'E�;8f�]� �C�O�֎��X��M�s+�!?���(*Æ'^q���"nb�b���� -D벎K��fj���U܅�b����7���Go!qΉ�*
�Y����k:�d7�0i�����ꌛV�2��~3�m�n-t��#��PA���Q$ #l��8�Ѯ�۾�B*%��D2���І�C/�J��f���f٥�]�V�c��LN`�9t�!��H$yo�*w��3��3�،��2H��h��'���;%�`n�֣�=`�D�)����ϥs�	~7�^���75-��?�y| Sp.�j��X�Ѽ��	qU�Q��A��l�4+��T�용�P+*/���XB]�8\�ZK�8��]��)�7�c�;I?7����-�e/is^���܌q�N|x������*�Z��隡�����q��%
T�2Ծ���ت2��������}��D��Fo�U`�0��j�X7�Lk5�B�¶X'�2j�ɘ������@�fA:q|�u����z���d���T�v�9���̽�d�;������c��p
���v_�ư�Iθ˙Cx��-;��Жl�x��B�#�;��C�$h�Ț��^�Nξ91JZ�g\IR��<K\	��kM�\��F���s˦ pG�~���Pt�T����q��?��Y¼mr&f�vc뽞�-�ڧPt0i�3i|����H�R�ྌ�Ħ�5$�<25o�(i�&�򴈧	��}���.�[�_�V
��������#�[����o����ax�p�n��`:HQ�R���+G3�r�S�1iab�d?oqj5���ßQ�x!Y���r�T�uծ����6���W�=�'�Ԕu��p~L�ތ$~�ɇ|4RE���:�0�#t��"�xy���#@��7[O�]Q��L<�]��v�2?O/��<!�MX�1i�O��=l�ޞ(8R3J��D� �b=�B\�#Ie���,���<5�cI	�\�I�,�����G�?r�����IƐ�ϓF 2;B-�uć�b�J�}ħ�E�6o|X����Ghy�_1�H�ČsjCI�:i�Os�k�����7�3���>� �����^^1�+����%���Te�V�N_vw�}:Ap��޳�V���WF?Q�#��=j��+:�Jy�̭�b+9q����&jO��jl��1%Zq�ٍP��DK��D�DG�c���1�P?�D`��H!ݞ���[�'l*ʷ���{R���-��ԓT����tK�&8��$��k(�7��nҜ���{����o�a�N�uճպ�Lg[�w
��X�}����T�k�4H�K�d������µP�D� l� bv-�5����~�^X��Д l��ە��/���
�&��ˏX��:�Q���č_+u�z��o?�����\O���m,��UE#�3)�_&��,񣒵���i�2o�kؙ'*�o!@�k�BJy��!����.mOA��72�c�(A�p�\��_iNr�A��B�l{���jf�涤'y	+��R:�='W�GlC�w���%���>�X��i�q紮���J����]��\�Խ�b���@5Sz#̴9'A(�%!aA͈�F��؝�dk��I�������Ӓ��m�3��)ܱ���?Yy��?�Y^��R
U�����Ȑ��81��I#|�c�V�3�Rs�h��#	)g�e����s �g�����F�
$�3p7!�#��VB}�q�3�6���[�)i�'�y�q�M���N~R�Xb�~�����{��Mo~̵���gT7�q��f/��.�h�2���8��"*���[u6�B�b�x��w��.3�=�!U���>M��h܈g!���@�<_��E�n��c2���I��X��}��Q~�H��w�ȵ>p͢���s��Q��v���?
?n����Sb�q@ax��VS��і,q'��p�����/	0��N |!G�v���J1�ٟt+�-~߭X�Q!�W��wB:�9c3�����'��?P�:��gT"���Ve�	%�[�0��X.T�e��\j���!@=��M_C�����nd��Ng�������5��q{�²auWW�߭�q���>����ԫo�L1���z��B��m�MI�<�z(Q�@��<�j��=�w�D�|>�]9��e�{;�n�3:߾`��%����>�C�^�����R���Ӟ�%���6��n"K�q��'r���x��.E��\j���U�)"_�p+���W +�r�{bA�G�i��o�ۥ��ii5+j��+���#\��J�
�TH�N�CiAx?�`����5�4GI�o���§��s
e�SH�LNP���y���!C�O������CywNv����\��翗��h�)ĞZe���\C7��P:�7��e�RK�⚏ϒC(��/p+uAYV�fB��of��k����Q.sv�
�@�*��^��h��P�� �\�5Z.^1S�AK.o�\\(E�S�~.�^�M�Z����H�4#�kL�E�Ď�Q:�90��Z��i�㖣�*��o�hp����	�
QOaWu�h�ˀ�ׄ��}�e�T�3�Q(&N �^�-uF�n��)ԡ77>R���au@X��R�K>�w0������|�}��Bw�*�q��3)��
���<Ǻnm�I� ����>�1��4x�����x�����փ`�t�V�H���=�����{����i��U��r�e��=AǺtc�4�T���O�ߡᙰ���� 6�(�5 �"Ξ~ЎE|n��̹f3Tܳ��ރi����H��`�S�V�+g�a��A��ƹT���I*�3���{�����`An���)��W)�c,�xC,���ͼ��cL�9�I�q���94
��%@ձ��@3�gJCC�B��I�{��u�ӗ�B��i,4.ܘ�륗QGf/�9ٕN)��9R���QD��؇A��գ�A�E^�ػ��8��+]��`���/�*��N3��ъ�]���`��;8Q)�Af�/��d*G>�R��H�hGEeoq�z��8���rC/+�C�&�������D�)�q�|*�~��k@��>i�X�b��l���vD������v`�~��R$Y#Q�����4\��(��4�"ע���[�����jW ټRU��b����Xfb?>�������꼍�c%�C'�;����+1Flxq8�&�X��z�L���G�p%�X|��#TSL��|��LL��	�^�5��r{�Q%X�MF)��q����{�Mݺ~�m��D?#��8&�r�/��FU�� U�U�)�������"ޞ��^kS�ش΍̲H������d=�t�#q���9���6�e�=3��¯��N}��5A7j��������N�wW�l 6g���u1��Wo�ڽO���CIK]ҍ4HȀ� C	ҝC	H7H���
CI7�!�����|ߵ^��?��>�������3�Ԕ�'L	)$L)$��uD���2i�};H.��h�{�-¡qזE��9І}s���H������I�E���F�����ل����Z�݋$��U(F��'u'�F�G^��������F(fHY#t��Ϝ�KM��K�b>��Ѿ~��"҂�Q���.1�L|�s����%��?�oUhŷ��a�u�މ�@/8E� `��\W�j|�gz ��;��²��0Ӎ&��#
�09h�ûTlAZ��ƞ��՚��;���Zws�>kӧX���?
�L�c��������#m~S�����7?�K!iERĚB!�V`�G:L�;ߨ�YX�N�����@� ��ݯ��jZ7O4:C����}ͭ�޻�왼T�g�J��E)�@�/p9��v�8����#y��� �c��v��U�l�ie�P)'La3OX���.tR��!7q�_�!��T}���vj�`%�[�y%��o�i�GZ���;�ՋA{��s�
B{z�_B�؎>�x�CEo����������0�����C��-΍�/�`dH�:R��'���06�
�ӿ���n��f���Ă�������7x���o���*p������t&b���-��#���щW/��OeTwy��rbF�1���:�@e��~Ar��q�󄡝�h�x�z@��\�'W�os��3ɰ��Z����^���Vboq���ǅ%�d�"O�>U��Q��#�4�%҇9^}�Yu��;��ld.E;��p\h�b��g�rbm�r���=�z�r��W���{�Z3a{Y��Y�B�t��P�H/���\;��9W�H�o�������t�� ���g��][���0��Ȳ���8��m<�� �=?ܤ��
�c��;�Cv�T�T�����_��=�-K~�,ugP��L�k3!]S�!�ޥjK��WH޺X��*5�J~v£�¿*@��+��Kһ�B��}�t�` �Dh4V�/�����{,�1GE`������"�IL�e��vPB� *��}阣��<�	.�?>բ�B�H�b�$Z$����J�Q�GX�*i i�;3�)M���K(�.d^��\�5WV&{��e��W��E��L}Et8z3��PX���;�<b�;���	�i�԰L��gPc3�G�Lt�{t������q�Z��B�/��Mw=v��9P������xP�[�x�)W�#i�j��LK�nU�]�ݦ�a�# sD�Q����w��e\刈?��vd�Ji4���y�E���NM�뛱�M��88n�dGLSY�7��7���j&��j�Q��/je'�Pq@Bu"h)�Cyy�����*�ي1�w���
�w�bhQ������g�Z�`I��O�?M�0f&S��Vxo��LX8���>����;*Z��7���
���,w��n����W�;�9
��/�>f�@����O7����ɿ�����m��ラ��.��Ł廎/M>�nf>��S�o�/ws�a͆�d<yl��P��:B��7~�U����5�
�*�Ѯ4<^Ut�e�4[�"1>�.��eq��~B��QM�����ԻƩ�w̹QP�j�U7#�X�:��5J����ނ�Uś�H��-Ax@�6��Y�)�,�!r4� x�y{٥dd6Ar;��)�z:����Ib-`�"��S�a{W�����̀:�Ռu$aa�Rq�0zX��7�K8�� �nȁ#��m��GY��{��N�]|�G*��\XZz�ʞ ��G9YeTѣE��(���g~Dӣs�9tR�
��uR�~�?��9:��vYb��2�������FU���K���ֺ�x�
DK)=ZI��.=}�����~�Ҵ	^H�X��`��9�3�-1���༭�1�X�Y<�y9L]x9n�
+��z�ˏ+���튛g��
�N'�3���x�cV7�dg����xv���j��gd>9FIT�L��ൻJi���P���!���ۖ����'��_Y�����I�^�s��H	��]&M8)3� 0��u��6���$Jl��bf
��_
�@��ˍ`G<�۹ń.|��]�����5紕�@���J)�6j"+j0�:! @W�F��|eh-��G[�܁e�rv�PT#�?	oP��uɔ����r8V���T-�f �b�$��E)���5\8>���ַh[�ff,�N��we�9�p#�qА�����|�C�C�*Φ��H��|�>�#�G�f�k+ ηt�i�q��E7|N0{\��[A��.���	�XL?�[ķ�v���W� �2�������˃l z �m���l�	���_�$9�M'��HC�EXRU�����~=#OA��)Q=CϱD�AT�GA�/�u�o�OH4�*�� ��LGJ�n@��	r��7^Z�pY"��2t3.�	Y�Y�GQ�����Cu���)�XjHhvky�,S�rr�̀�+�S+��?���5�}����v	�&��#�s�8J����=p�4�� Y��X���n ��:2����� �:���ӥ+'G�<+V/S5!q	�ؤ��a:s� ��|��p�0g���� =k_�#qF?3��DJ*W�z,��r�k����!� D��#b����qq_bWH�uװ��p"ї���M��L@$��tDa��!Y�A_�r]��3}XW��mXjB�;�
�U�;�ߠ��O�Tt���d<5b"��DQWStr��\$7~k��',���pU��)�X ��.� 3!���d�������H�na���F�
���� AP�z�#NF���h1/Z�j��:�A��w�u!�������1xm�ޙz���#3)�?[������/��@W �Ik;4�E������
�sU�v����U�e>D��n��2'����"~��H'�_�e���3�)��>c �<���Ǽ�c��AE��+�$���c֤pP�]x��]���u��%�b�����dj�m�}\����0��08�����_"[Ym��T)����[s��B�o�q��A�I���L��h�>:���LR�̈́֒C VS34fT���J�v����g�bix���F%���A~V}��"n].-�ޕ3��~.Zp]�R
R D(b���~�jJ1s;��"��*#��Ik�숎���JW�N[0��߽{�Qj;��j�ZLi��rKy����zс���G�L tޟDp��x\l�/�Q$x;��׻�-�p2��{��6�0�խ?;�#!���g�1EX�a-�y��`:o�P���6��"<.��ޛ(z�w��eZ6��C@V%��ۍO�gO"8Q��Ln� v����-�������+!���-R1C���>^FQ	�t,]Rٌ�l����NW���T�]$_�������<��ӊT�Tj�	��L����Ua���p�ꀩx6�-��:3'���WŪ�1������8}@�6�籜�j?9
�w���o�]���ś�eSF�qI�0��]���ľ!c�i�sE�ԟ�ʊ�g郬f5Z��v8]�!���c�k㏇)��u3��mU"b������ �t�<=Q�ʈa}�:W,�N#�
Ç�srh�������BqI��������}.���g/�1
�fׄ�up��c��]'n�AN�/��72�EZP�a�����-�-�� ޷F�=�*��f���[�4��g�.��:��.���N��E�3K�yx��Y�Q�7�FN[�َiϣ�$a�Pj[��
��9� i� �=M���:E��X�K�Ǭ��]�<��zj�Y�(jW��������J� �vq��Μ���1YW���V7���ه�ynR�зB
"���J� �Z�Kp�0~-�u�.��ʏ���Kѵ�A{�����$>T?�U�"��,�%)-�6���ғ0$!.;���D�j�bl�2��?�pA�@}����˂�_��#�0����_����L�?9�ʝ���|�_GZ����j�Η{҇��0`��N��S�r3sldG����e ��w`�&B��F��=�\Mg0��d������[�+R���� �P��)�'�	��!�S�����+O���:ztY��;x�K�ޭ"���͍kB�CK���I�f��9�RBem*�3�Ӹm���wW��s��H!�U�G[N��3��# ��`�r&�o����/�cl{�$�����=�K;�y����/E���
��tC/J޲.<!�ο")�ep\�~�$�	�~n}��ďL�XI��C�:!� �%r��:n�%1��|�8�^Cђi@%��ˤ�:�;�3~�3*��������|��߉������*Q��T�1��Ź�r�� ����v�L��(���P��3M	���S8�^$��|,Z�+�g�X��P\l����0;a�z�i�g����"*�m�o�a�oJQ�d���Ȯ����������Ӛ�U���N&�;�j��}Ō�[|��/J=���M� ��L�~���U"ѽ�JR��PiQ�'0��N`�Ԕr�^"
�b2vՖ�D/�)��X_A[EQ�YP��7=��\1笆��$�<�H�`��7�bD��xӣ�7�����ba @l��
B�'��+T�Tʈ���Q}�H�ܿT�q�=���ba}���94'#B�{�#�+�)��M'h����䠷�a��^��=���)��m�QL�A�v�Z��!OJ��%�PU>U������T�nQL���^��,`�Fց��>�\�Q��y�B�/<��1X���]�Y��C�st*}9��ڧk����ߐ��w=Mbv�g/C�}Mǻ_;�6�cm̬�W;��:,?�4��Z	$�KV�����_��p�~�-#o ����=i:�mT4{�s����t_�g3���J����=��D���t�1�'��@j����o�d�qS��%�H.[�F��:b���z4�1������`��K˙��OL��"��T� ��ͥ���2
(/�a�{ݞ��&x)��^�1 >\�I�����w������~�� a�0|H�)�Y|@D���m�w�r���t��a9�>�@<z�������!�h���Q�J���tl�*�z�I��E(��j0	�
��` 1}3������o^5��x~e
͝n�v�6��7�x���GB�T�}'_��Xo�}�t2�<q����i��'�I�`��Rၳfj�@��*�I)+�&�1����=�_�M�m�T��d&H�*���)^��e�8{jP��џ���I!��N���srt
ݳb��~Z�$��?TnU�
�NƔI$G߮~3v��Nmt��γ�Mb��T��}\
��0IđO�]�|�W����e5�
9�l��3���e��~l�)3�1\��q��ƹ;}&��� P�f�� ��jxۙ�bV�D�s�:2�k�g]�ų-F��ު@�kה�|��p�Mk8my���b���qm�$����ggS�M���_��\ԅZ"n��3#��9���)r��H���/b��
p �^�=�D�N+�X0~A��5��T�NnV�}$]��Dq�G.̉G.�JF&����-[�e+[��|磖KY����Ӊ����G��o
t�|t7Qr�q^~�u�[[�*�!��o=�ߙ��W��d��^[�%�����a~A���uS�V�	6Fy��Q�i/�T&���!q>�8,[*hE�/q]
��&+uFx��>�qv���4┧^#�w?+l�$���e�4.�.}�aTnG����Y�R!���<�-�
J4��{>J����P��;��@�Q�)�]@�� ��/9�ҢNh'�I��i2���t����N�p$�У�Q��8V1�Vp��e�N�~�J�~`�?�L��e ��)�+M �^� �g�/�y�:�3E~�N�)"e��V0ė�[���I�\�.D<�?\�����>�������۹s�0ѯ�7��Lg���b{�������	��_-/���R��>}��W�#�u�g�H�l�&�`:�}��|׶��ɍ?h�n���0R�9n��d�1�z�����%�P=>f.!���N�<�Fy;�	~�R;�����nx9�n�̷mGo):2�*�
T��N�x��Z��ϯo~РU	XE��ys�yzydN��U7�I�wT��3�ʑ��U8 �4�����Va�t0,��E5ՆfL�LH�I	݃S@5��:�ɦ�*LM����;J�w����n�p_H�$�&��R`�b?�����8��R�{j5�T���a��/l,b�� 2���Eџ���j\tEo�����_/��(�����KJ9obC���5��Gi�fd��59�>O��/�L��2o**׈�L�+�����<V�czRs��^gH���,a7E����n��Ӡf5)�`��4�����.<�sf��Ę��(v��6z��F���_����;�+G)ݗ@�R����L�ˇu�/h�把T��j �e�w���Jo1�c,�'&}i�7{닏 RYW�A�1�zGN��]V ��piٔ�▴]�����1���r(~ݟ@G���?W^���"�����	�M���A.�䙸 ��	�8�o�Y��o�4ӊՃ�>"S' \���ͭ�!@�!��C�6�-o�_.��v�5m����<mb2�Z����8����K�2;.%Θ�:1s_IM49�k����z��]�4R&�����NA���>�DF�s��Y�( 6b_� ~\ϼ�=�X�©�}a0q��R�S���e���Z\80(��çFo�q���Ʃ�/A}��:^t�����B.�Z����� �f�s�@Z*\p���m*�v�����g?�1
�T�;%���2?2TL�G�H-����윲�KÃĂ�TzK#����K�؅���CWp.�F����:3tg��'b"E.���	Im��ؿ��7=�i����-sk��u>�P>!ksO��^�����2D��|@B�<L��v�{��[�5���'�ִ�*��=�������r>k��Jp.:�}��휦I��%�ڗ`N&���͕��ez�YB����	2���������X��*�vA���y�����5~.��އm$�U���
��HYʱ��R ?/w��L�����]�&vT�����X9�ֽKL�/�]$�gn� z*H��4��-���?L'�K���P��^�'\�?�>����	R>�|.<wE�I��C@T�4�(CQ�Fᴤj�����XFС{$)�r��o��R,�&���� R�M��(n��ϔ�f��txQ�D�Pz�G� �G���b%�ٿN+l`�)�Wwل��6��8�C�[(�B�j��}�3���l�F���!O��Xޡ(���kb��V+ҏc�ЋI�7Z�}��B�&��n��R���ݐ�5�k����MSM�29e�4�͓m�E�E��/��w�	�^حUi���Üi��i�d���
�p���j��l�)�MȾ��a�B�u5�A�����s����i�z������ڝe����8n�3������@ɟ�>��F���ZuE[{��M�n��w���E��G���Y�|>���ґ��QN4��'��4��gR��q�3�PJD��K��BG1м���9��C��/�ʭ5��G˘����#���$�KA3DP]?�����
X+�f��'
P-�>)��Y��(�D�Y�^�a���r�@�3�KҶ�A�hW�j�)c��a�5�u�<}��lx
���ViP(�y��wx��_?j�P�9l� ����?�k��7+Ӎ���3c�+Dj;�-��'[����c׽��Z�Gj��l]���X4�����GE�Sh�E���?G�]qs�2R:���� Ռ�x�'��X��k,E� ��ih�֟�9Ӷ5��&pqN��O8ޞ��UhU�0���s�=xiE��pM�����n[����F���.!���M� ����s=�'tt�2,ir���ؿ$U�X�N�~�������C`�,��>&��z��4�'�
i.�K4{�ha����)'&CJ�8	�N\Gq��Sh0Ć���>q�������ߺCs��E��
����Y[�]�BQ�K_��5&2T�d	V�#�$�b���w�ϯ���ᰶ�N��K����r�Ҟ����"�5,�/6A>�>�o,Y߸QR��D�~iQ�(
e"�k̈́�z��
5�L�1�P��c۫b�2��f��y`��=b��^��^T���&&�,�_�:��� `#p�#Kd�����ϸ#]Y��١Gk�|:>3s���4v���P� "2��w�I�ӯa���u?
��\�y~cy���J�@�V~l�Xt�E��G'X����+]� b|,f�����V��9%:'� كq`�Y�qA
�9�>� �#x���C��M5���a��	8���<|��S%���)Ǝ9AA���nH� ��o
w�����)��m���,�S����Rw]��$����~Kv�qk;ߑ�m�8�֓�;��$q�����V5,e�n��H*��VSF@/��Q��*CE�����/�s��P��ź�c��l`���d~b�O��Xl%�����Ŕ���V�����5��v���T��gKD��#�۠�?ե�V�='�7 ����@��ԑI:��Q���m�So�L������!G2M��ݿ�P����sq�����f�2�]fO�ғ���<As��\�����sv����h��jT��*+��F�A��P;�[���=�P����;![eG�1Jm*0E�P���Y|G2i� \����ַK�6�5�փ�Xlk'��?�o�+���jj"3�3Z������a��(sG���79��A��rzY� :�T�Q2ϫט`(
���?
;�>ջ�>��k=8�b�<��*9Y��{�_e���X��TG�N��NW�4E��aS۠E���G��V�6U\�Ys+�� �I�s����?����V>�2�D�>L������<)[$S|z�,����g�_�d�1������*�~����zD.�~.�h���X���UJ�d�USi�u�P�d�P�I�4S�~��R�ѰV����խ��ȭ��PG$nD�'�b�i*:NU�(^��)k�L�b۳�����)�xT������L)ɠG�è�_�J&������z��i��\QErn	���h�4͝���C�4�	�V�f5R���J@B��-�����C�&��?�<�Ш���* �g�]���["���=���&��?a����h�F���vǭ�L�\y�F��ΑC�Nq���� �����E�Q�C�"�)y�qS�R���h6�Q�	?�XJ�v�t��7!�n�1�MN��_C._��lnN�9W'���G�ۍ������Ɛ^#�B�
!N�ܟ�+*�T��W���[�*���+G���W��5:g�˅��]�������~U[$p�+�)�l�V���.�y�++l9�&C��Ľ{m�c����|�xŸ{�
e&�F�U��#���DW-��i�9��������u���?X!hƋ=F~A�G���-�bl�>9\Z
b���@��#���Z�ll�]�1f�����{�|����~u�w��������&jK��Qy���d��2���˃�������ꖿj9GG��<���Y�����[���Zq��A���FCՉ�JK�;9�O׎ּ�OEã	;{�m�W���~��	ͣ�<�$R�)�^��4*��?;m��i{>�$�5�6�18T�Lq�V�@KO�{��;GҫR��G���7�	������{F� ��>�vs/���Rσ ���dve�΢�tL������� Tj���J�̷��]O�D�¥�X:�3�G��~�`�4�В���B�A�[�����&���kI�b�cu��I��)�|����M�^��
�/�,��ܻ$*Z@���g���:����I߲�8�孭_
~m����O生m��>����_���o��ء_�Y�*
�Yer��h8���q�c{�����]RF��·���tO�x��7v塑/ȿ6���x���O-�p�T�YT󄯊��Ô����lu�{��M���ʙǩχy5��>4x����I3��'��(T�h%mI-�����a�Se�j`�@zcXb)��4C�Vb�Z�.~���)�Y���ն+ҫ'�=���� ����� �_�O/�ׅ�bX����KZ�3mm&�Ֆ�Ei�mH�]�	O�)��`��������5��;9�D�ݣP�$�ovin�u*j��=eB9�)?�tK��Z�P�b@f�e��ߓm�k} g~��/�+wu<yt�=:꧝��V^��{���l�Z��ȶ���Of�os���h5T$�T�@�*)_r4/�2��G����d��z_���f?7�Qz)������H���P�6�l�J~�|�g����-Y5�)�ܰ6*����f������ ���]�1Ϝ8S%�J�g�x�;Z�_#>��sC�ZK��s���i�C[�ţ�u(Z	�˚i ���')fU�9��B =�ƂiY.z$S�G�<�F�Nrx
��E9 ���r.�a>!\Υ'U����}-b)Χ(z��<��|���.��X��V�L��JŁX���o%b[��k�/GI-�f�ũ2<v*Y����z.��v6�+�U|��w�]����6:�͡ܦ�}F�$rg�L�_��P��a�H	H��� �GZ+K;M��q,ǐ�z��]s#{P��at�yt��v=N����ku��l�W�C����	�"f�N%MT�P��&~�V�'{a7O����3������+߭# ~��[Yϊ�Bo0��PM�QK:0|p��c3 �D�II��\��s��2�/�W�c�Rxo(�$4�A�s<vx�Gz/��_�-/]ZVV����oHl+�C�~[�r��>1�S:R�G��1@�@�7��p�/%�z���ӥ"�Ș��d���ݵ���.�x�l[������D���%C=ٓu��ʁ���+~����+�4�$J�䛲���MpӍ��:|Xʿ�t)�0�:M����l9���-��sW�����V�c@K����RX;�d���KɟvBs �`�.��8 n�@���ZyT�J�-�P=�/ӿ6�0Y�球aݻ�5�=��AD��?��ݟ�i<�_TNo~���tB�}"K�����]�!)��B�,�(�n�5�}�Ζ`çx$��4��� �/@_�C|Q`]a�ҋ��{m;��]
��|��hI9Yo��E�����m^�r�+WO�|����Ǜ��=_pl>��@�?�fv����S���Y>�T>��+h�փ$�uYҔ�T�+~�3)ǹޒ�I���>P��B�j"��Z��næ�S�_��t� `5�"���V� �#b/��{�P7�A�,��P��z�*kbA��28�ok�YT��Ъ�a�z�o�/pcف��Á! ����������u���Q����g�?$�7��0b��ΫƦ[�?�I �>[K>��֪w��%S��%ܻ8�������&�q����X-�w�2U���`���n�����Җ8��R}v���uK���`�a5c���?Jb���@��O������v@l8�r�"  ��P�EQ�81!�+�>�l���"e�����A�z�G��:ݧ�P�c�y���zǇ���þ�5xE,�3Q����A7��o�������;P��7iz=lG���ޝ��,m!�C�^|2��r�� !��e@���m��U<0���m�ªb�D�K�����֠�ۀ���/'��t?���d�G[w��>K�bN�y�*lG�@��eCC�Aʄ���ϡ*�pQu��>*wU�(����Q0x ����a�Ԛ���X�q�"����,XRi7'$���`!��@��]��TKeIA��`9��r���"�We�h�]�T?z��X:���v�cI�<\ё1�M#�8�$�t��Ǒ��^�xz�s��cqE�{{u�a~�	�fK�R�L#o�@�o���'F&��3���v/��-���۝=�%���S;�>7����OV�P���5/��SȮҜ`���:-x9�@�^�x�2��2� hGi�Z ��l�v�2���	�z����?w��#�ۣ���9��+����P4謊3���ߤ�ۜ�'~���%_�B#�N'ҀN>�������b&�Y`d�8��9-�o�v����j����(�Ex�R��p	��Pϒ,L�B;k���0���iSx�<�S���C-^��\T�]��0) �ۗZ�e=˰+�����b>QϞ�Pщv/3��j���dN�x���ux��ǵ:PK�S1>���I�n��_k���o�����w�ѱ���:�b���,�����[���8x�vƭn:h(G(��:}���8X���T�ہ�@�S���̍�7(nN���r^Z��bN�5�?U(��ҋ�A{�[�7�a��?�n�6(e���c+4z���Ta�[]]͇|t_QrP&\��S��;mr}�u�I(�W������I��A@k͕_�mA�f FG�Y�H�K�=�E��C���bٺ"S��!I�<mՄ+g��819�������R�ա0	n��ovK����ͅ��"��1�{�F�%:�xg� °��eW�M^!M߄��?b#����zRDSϞ�ED�NOH���D+��{�?��Wۯ�\��%��2+�0l0����p�߀�S�v:�M���~q:���n����[����ھ,�'�N,{\�s����)�B�L%��-/1:K�&�d/�us�E59� �W;�;E��FD���=������U}�)a��pR���_�����Ş��B�Bf�y�0��4`~@9��0b���̂Kv�8��-3��3K�Q8��pS���歴UC}GeOe�.�Fk�o_ϝa��-�~[�����\�m_�w�,���@S���.�P�":�:!��L����U��Nw����&Ɓ�jX�uTB�#�(*ml�	̄�T��VG a�g� ���{j$�Ӏi���S�� ��x��߅:ح�}c��1V���E��v�w�Ɂ���1�L�P�ϣ��GӣQ�� �th#oVӡ��"��<[��^`��g}�/�a�_�y9��=E��t�#Po+�ZC�tP|���U��);�H���_}X9�>2��J�:�ͬb;�HN?�%J��KbW��s�ֽ�UQסZ�R�����V�)�Ѱ�xuQa��|�Y�V˥E��9�b��)<�O��$�@�bL����������&.�Y�t(U}�� ��̲� ��'��7�����S�#	A�
j�a����	-��s�;$g�3�M����֠S��w�X���y:(�~��}�t�BT�v璡����³_�(�;���҅��I-M� Yh |�4г�)�f��5�v�E�J��~�p�;��PblD`�k�Xl&sQ�yO��~'�.گ[ � R��v��}�P8x�O�ao ���	�]�I�=��l��yU��=�q�!��'�w�cH�B=62�H7J�[��2�A���^8Xl��4����ɣ�"�,���䍮t��}��) ���L
Ƶ���ߠ�Cx�l	3�ߕ���'^��	の�
1TY���Ǿ't	�H���Z{�|cUF&Ӂ����!M��z�ik�	۩�wbY�b&��.iC��B#!0�N���c����?��3�n-u����î/�=��zJ)8ue���փ�ޛoXf�	۾գ�/^�)����M����O�P�3�*�]j��~�Q������~�(X�UX�zi
T�V,b���DagC+����@q%��z�p�AU,qE�?�}�M���/��8���/��x\�~��n�0�
����+U�,g��v�c��-V��uYDA10>b#bW��{� టs㶒3�����#�֛��[n��W��R����V��AMK�S��rR��^��?��7z��2�.טl ��sy�g�k�6%GI���`a��ph�v�D]y�AQ^�ڔI��!�7 ���^��3�,h���D(���0�:����� AQw����nR; �gÎ�^>ģ�����Gԅ2ɡQ>�2�������AnL�#H#�C0�
KY�M�&�;t��]��.;�L�1�b�Q���~�a����w�Br�!��l�kT2ϒ�����Š�ox�X�02=�BЉ��.��H�pM�T����*QɎxd�n��}
� ��P�bʾ\:TL(���,����(X�%�Ǧp�:�;Q��A���HgZ¾
L+��%-;��K�u�ȏ�c��x��cY<�e�z>�qNC��^����`Ș(�:}f,<�1�sl���сԄ
����n�K���ް��X���*:�)�4j!�ЩP�P`LL3��+�F������w����osδ���5`I\	 ��o��Dѡ_{acg��8�����
'j�.�Hm�1կ$[�O� "�D�����n_���䇴cg=3i��DM�Z �|�ZKɊF� �
���]�!:7�{��9�t�ɯ)�׀������E~^e	P��H������G�unp�fޭ�����n����D�U�����eQ�^	���J/�#]�󣈓����Q9^��F70��"�8�&q�%̯�ɠRx�X��_��LD�;kEmj��I (���q�6TOwD�3`�oo�G�;6���M.��<��=��@ ��q��~�o��Z�u����۰q���F+����FR��k	o}�F��>y�U�y2ۓ�1���θ�M��j[_,��\%�E�D�tˎѼ�L�=�h��L���k�M�1;�ʎ|�.'$���B���5#t�U�sv�h����h�mj�FdEݸ�><JC�N��
Q��xq��P��"�cj�bb�f�=In��2�|�U{�s���]�����omwrF�x�t�Z��t�-��R~@��J�H#ȼÝ�p�<-t���6��)`z��v���=N�@�zd�=�@#���ȣ{�2o��*����X�UY^��!��?k\)a�1���*� /��Y-R����a�p�J�a���j��Vt�������`�+�ե�Vj2Xiz�����ݨbV�����[8?Mks(d�v��
	ޏ!���M�P���T���� 
0�R�IN��I��	�b� Mo��\`�>�F>#/�XU�]H��k&�~{�l涖�P�Ǫ вQm�8 �PF*�Cs���竡�s)A��ݳ�h�����s�r�B��9�'_^�>�#��hi|2���#��������t햑����8u"�{����tzWi~�c����c�_|�EiR�}� ��J���+f��ں빤����,Uls�p��C3-f{�?��(�����]q<�B�����n������!L��% X��1fUJ����PЛ���L]�������xџ� �(�|�|+��q)��{x��+]�U�t7.��	�r*{f�'YCi"A��D>�g*n�p�\[]�-m��Zx���Wĭ�����?�j��'G�<��>��L��k����[��b/�|,��H)��8�0v�"E�@�:��αDы�<�p��۷8UƼ��[\J>sx鼅&�8\�ѧ�̻�u�W8�G�p".K�uv�	h����Qx�F����_W;���%���?*�?�ai�	���L"--�����"-C�h݋����9!���I����-V�NFpk�����5�b���y�InkJ:�Na�r�GD܆�V��s���5�+1LI�;�[�ǤMf���w��D�_d�iob�ӆ���KV��T��T�+s���<5��k|��:g< U{�Y�<͠�[��b��\�9�T�޳f�'�j��~H$zw�,B=�5X����5M��9ƃz�<�Ӫ�f��߶��WZ�|�8k���Ky1��[�<����O"h���\z���*��y�ޯ{���!�G�7=B�v,ǰgI5�|�(�42��K�=s���)L88f�^�`@@+XE8`������bi�U�{ѩkև叽݂����V�@80?{�O@¥��������g���},k���(O��=��7>���kR|4V���v��W'u<	�
9���z|�S�a����ص��m�UF�FXW�}zD���v}t�fc�������<25�߻?��2����ϗ3�#�k6o� ƪ?��.߳����R�<ׇ���*��#�ȡ�bU�)v^#d5-'����ק�qp5��\�k��!+�(s��AY)��g k�.c�sCt���$A@�u���v�ȣ���g��[V.I.�Fe��Y�̥���6��H���9�qqd��gBx;�ٔ�m诨�qw�}�)2�Ðgݧ��Tj[�|���h��H��$y�Έlbor�w�x�Zlv�æ���pH����NK,�u8�5� |W�r<� ���/�eߛ��g��$2�4*<Tl۴G����ΛCiKF�U�8�b=�fkm��U��.���#�jW�'܌�ZJ���뢏�n.lg�i7=��,h&=G�k���C�*kn�
4�@�R���ܫ��h�NJQ'SVS(�U���o�T)_-�o/�x���F���3��c$���6z�3hS�k��H�L�9U�+u�8� ����|�$f�����=�.~�����
�i�2H���6�Jb�n��ȤeFr���*�N�Ft\�2u'���c��~���Q���9ݍJ� �I)��!)�[�%�C���
���tIw���y�<����^��}��}�u����R�L�떓Ō���a�)%�:@��8!#(���G�b�DN�/uD�����$	�B���6X!��a��`@��6I�0r��v��t��T���3[TW�u7Aqޕ6�����,u"��D�Ԅ.�q-�/������8��?��z���^�=_&��:Y�����~@����}���==g�=���,*�[���5�H+H��|,�S�8���3D���vh��gA�[V�����(����y����>�:h���K��h�!��#����5$���ݯ�
�����/��(	�+�u��pb�o��^�X"����.~�l�;"�sR�J������p:G���j�D|F`�"S�l��+xO�`�>�_��O1�	]�B}�U��d�U2����{]~E��N�� �e/s���*S7�?ڦb/�unXo��r��k�V���+��~9O��P�w;�'�������p��8�%�$4|��K:C={�@9���{��a��O�&=w�L:}C����
W��w�qwW�B֧�2��n�>��uϯ����RI��,�g��f��$�"�
Q��Ð�,K�(j�4��+}��WY�����i���撪J��{����Xfz��(չ�ȳi�p(�kjϒ<~d"i=6w�Q�7�
�+"���|PN�������^|p���mM�+P@N����~���]���<n'P�On5�n���qZ"��'��m��5��(�-� ��9H�BIѲ��G^/�d�	��#������$㌥ִGb:�Ōx�Fq���������@H���f���Duh�jܹFօo4���}�}7�}ޥA�������>K�$�ƹh���j�/J����Ka7�ѧ|�1�Ą�!@S�1�ə����d���owߟ�*�5�
Yf.P��OL,�����jI����D8C�>~�ĕ�D2��+K�r5V�m6o�[H�/��r�;�l�6^��� ��O8�H�	9���{Q��ν5����>֣&�n�,)��p�Ɓ���L��K��#�6ħ
�ɗ�ː��d@��!�R	����^X��R�Rߡ�*|@!�e�r��?0��'���e|}n�4*� �z�3�y������s��6��<[g`�w"�5�a�_ -��2��$�G�g��EP�~M�̲��sY��O1����B�S�l ��̡�?M6ҏu�oם�R�')G���œPP�"e�:���*,��}�vm�r>y+0a�͐{���O1�vH�^Y�f����N�w��_IL*���Ҡ)��	�ҭ y7��f9��6�CZ�C"?mq��nas�1���Z��gP�Q-獼ʌI�2��RnTjk���?�B<����o�X�����3�%��v����V�B�y_Y��"2��S�m	
}��j�z�EX]��{XԐmK$�qW�G�n"
��t��̋�}u����V���L��J�mB�n�4�}����?@����Z��zɓ�$��; �ǻ�I��\k3�R�su�惝$�:��>itc�T��~����Y8�ǁ(+8��ut�U��ߒ����72��q�dƅ��^�Upy�z�/a�A�?GϗӠ��hY��o2�&[|$��K����4,/�J��1N:�D�ɓ6�2�l�$:lh��`�._��-�θ\�Ml�N�s���($]�)��g����z����k�a�c�D�O�q��ZS��E�{c�'j�h�!˂�����r����uOjizY���+1r��'�w��������	YX��E�:�vv��??��_�/M�_pOآf���;�O↔v��ء{�@������2U�s�+$�v���뮜��/	�QO�[��>ƿ���4�:&�c�ן&D��҈}J����G/��Qi���=�-��v�b2�Vi��K�5�"h��� `���
id{��9;�\˵����0����W��=�H��&4���Ғs�M�}4n�N|�����O�B��,Ug��8�v �r7�1�0/��,2��w=��?mY�:T�$���'�	��}���v;�p�'���W��� ��_��-�z��s`u�~~���v��T�|/�}Kē�ؓ���^���1��u�#�M��c+>�c�Fy=k��\g�1��I��A��O�[�;A^�K&�z ��^���@]Z���{\��헴�(��8]��/y�/y9���x���'�+T!��:pFji*x;f��	�ځ��l޼]����%�h����/8���:�|8?��V�+ #�J�%F Y -?*Q�'��䅧�@�{�:�s��ax���xT
Ps��]��{�)��Ѩ����@��wֶ���i�D���}!R�ͯ��⤸�7x���e��B��H�_����΂� ���@_���|js�ɳ5w |+�t��K�~r����.��ڭ=ۭ��j�X0LԷ`�Y^_�A�,�M��Au���`��޳G3��M��˯g�G�gxIW�RxOtSJ�d�?~܁�����z6�L���ઓ�\G�3E =#��i$��,�<��
nsE��ʫ=��+8D0��[@m.
���ğ�08a�G��x�X��P*-��J1xn߻�(��D��C�)f�5��4�cG��A��掖ma� j|U��]B�|��N:��ý���/8���2�޸c6�o�B?\�⩽ZC��n!�Sz���v�w�o��87����/����W���S)���ޝ�ȃ�]1镍�@F�����9~��N��~H�!��(���U�g�)Ak�,���I��8s�c�=G3NDUy�2%��#~_n"�\��=���A���y�h/���<�v��)��]jҦ�
s=TW��̙3�3��������3���Wėi��@��� Z���ԩ�D��,d[ܶD���7�W�>�������_��?����enz��A���L�;�QP�H0:Wrv�|�u����/y ����a�n�~�+�㜰
�*ʹ���g˨W��̤Pvq�B׹֫Ƶ�5�?s�T�I���dN�vq {��n:p@���P.�ɞ���tsy0�5.]�jC-Q����e��F���_N�'�"!n����|�>Z,��q4,c�T14�?m�����"�}��i�XJ�qv���՜Hu ���/�p<�D�bLot�<�F��o�
�! ���/�g����ajJkU1W��K�s�QAF��Lv��]�D�O�k�i�������dZ��n`eaEj7�(��X���
_es�bi <&nR@�͜/��i"�	�@�h��~�e?�6*��g�*'����8�-s�8+�a%����JQ�oƯ�d{eܙ�I���V�uNZ�{�����}Ń}�[y,�&2�@��-�\a��F��,��yʸK}pq�����L�{���w�ޭ`,�r��,��u��^��{�r��u�.�DEQ���r���Q8pIe%2��"*1Q���b�_è^�p<�R�ӫb�3��'�<�Ӏ>��܅O?��):�YT��L�m5�f=�T�
���s�&������j�z������alˢ��J���O0�˨���~:��T~�����h A����n�o�Pͽ�5߄��/��o^�֎�`-0D�LR�
N��8I���KV�?�Yj��JD.�)�[���)A��/��7
��3��Ơ.�N�z��;�!�|�jo�9�5X�q������c�щJs�2-�
�.�c[*6	�Ƴ�E1��4��1"#�rløaw�y�Յ�4�	����n(���\��x�a���KNQ��8N�{ L+�9��0���+t�i,�6G22=���%�i!*/ƒ�Ø���a�A6 �tO��e��HG��Ab�(~��8��V�G�5��fD�x�]�{���#�7o��� 
� b�(�A�/بPFe�7��X���0�Đ�	GtU&�'��k����W�1��O���v���V�'��W�[?�gL{��{�a�%�h�Ff�bE�Bc-�@���ܖm�S)���\7�;�}=�X^~�b�-=�����CϨ7S��^k���������uH)]���èxWS��
���T�꺴�z��w#�&�dm0��� ���œ�lONx��A�<���꤮�y>�Ğ�O-+ͳ![sH���x�E��V}N[�u�����S�*׹D�|� =��t/��=�����m�%� ��}\\��<|�� �!�� b{��'1߸��++��P�ϒ�/y�W8LgӲ��&St��c�q�����$�[m���Lk!j@4-aNT�jE$����d�����2f��c�,���7�s���8�r!k�k~D�����D8���O�w�
u�U�Hi�/�8�D~����t&?����t�z�Ħ��Ъ��$.��g�pD��wI4n�]��L�f�$�� �V�?!f����o���Yz��9� 冈��py�@j���$��HO�U�)��u�ܕw,$��z"AR����\/X�!Tk}�p'`�c}�b����<d���z�yr�!��B&����}e����f%�4���u��j{
R�̂�%r����>�GTbFq�)�xX?��}��\���}n-�fN��ɌHmEJR�vel��^�j����\���}���Bg�QCg��N���ޗ����7A�Q�2`�2�c�9�\�/�.������m|��]��$L�Յ�_Mꬄj�V*���B�����'��|
���"�����Xo����q[�Ax��o�_%~�n�G~(d�$��L�+�Ui�"�G�������w���Jw��~��&�BD��eU�Yvd`�ho
;!Z՞��2n�k(�}��jB)-��\�	�	R���/O�CI�������I��]��&��ǁ�?���	"�����+�����
�x��$�S�[VT���Q������� ��Ӂ?�B2��4]��)_%�X�"M�U�>Zp8�<��0�N�Cu�3���	Ӥ�&�@����N�E!OϮ`�{��R�ԙ�'�@�wp~����r�O�����I������g����fxe�a��ӡ�3����J��|�>�V|ĩA�1��B�~���cDW�]ƞ�{�a��\��w��&ô�,*N&�|ʫ�xHu��态�OH�*���_�|�7ʪ�U��z"Q�s͔x\D����H�=�&z������C����饩�赼��u�+�,�ݗ��X�V�z��~Zc��X>�ƌ�]������L��բ�B�ײpY�[��l3L��B�;�C�I�!��
0���N��Z�uގ�g���}��*��"@M�L�ػ�$y�i���£A�!�QO7HG�ڞ�V�>��"	������ױ��0;��Z��l!I�pG��Ä��qw���Xoo2ra��{����w��X��P��/�f�d�޶@ﴜ��ҫ�(���ߢ��Ǭ�4��(<\�A��[㷤LҲ���_�-"�H��TY�z�x�1��>ȗX�,�u�������ЂX�PN���7�{��܆���vg�\���s�*vqh�W����Z��֭4��璊�6i]��S���[H�u�>�ǱZ�Z���?l5i>ۆ;���n��$�L5@7܂'�䜔 Go6\��>|��,��YA������tM��PWS+;� �B86eW�\�:	|%AX��*4���K�j|b�(RFp�>k��x-4�[G/C����������z>N�gl�����V"�q��&޹��+~;�:��CĬQ�~ڭ7�y1-_e?Q��"����}��fhzT'{��d���2�D����t����CƊ���:1z��}*��@G�o�r��0�W|͔��f
rHkq���=s"�m����Ƅ�����(���S��g�l�Z��N���V��Ȣ��n�6�\�Ry�d�:�ŜxY�s��L�����[b�З��z�_|�G�.�F�ی?�~1���|�q	nw��EK<8��|/K�A�ŦR�E�3���rAe꣇�Ia�u)�o��������Kb_��ߗ�1�=<�p�|���!:������
XB�8�I�d��D���i$��/L�&��a���~"!�DE��nw��1�u�>T����qU����ԝ֋� �b{�<]«@U5���?�A&#�^�o��j/'��6빗䘒�1:fl!qd�Sӊ���MH��e�k��+2zR� � �r%�~APi�D:�T�;���M�/�U� ���er:4���h�+qx�����Bo���K[�^DFeڨ��/烒ڴ�*n��]@Z����k$-{�f���d��.�PY�*�&zb��׎��8�%��);��!'q�8"1������n�{�C9-�@9��d�I�������P5FO,�t��l0���-���Y�C�+�m�N}@]��W��:ƚ�A���k?���|����k���#CHT@Iˁ�N"�B�G�`Z��33���BEy��c�n�7W�����̠��F�����AG��c�OZ�>���O�k�oޖx�`�4_\x�]�G����±�n�1 ����ɱN�rw՟#��5e�5�0���
���A�o	���.to$�:�*�_v��Bfճ�xh�N?���8M1�5|�=��rҥl	0F�+�\)��0�.��D���~�&��/��*��.�s���Ă���<a��p�f�NJ�$����s,a	��+K��n���/I�� ���lW��~�-����ۺ����~S]k�n�3c��ń�E� {�e�E������^:�F�����f���0�⋁n~2���}iC�|�k4�t�5[b}�ߑ��%��`����UĐR� �l��_Ot"��������fH�U$->	=�7Jj<1��"CHI#G1��֖?-�_�g��H
�Kc2Ti��%HQ�:��0} n�����G�ŀ��}����*Q7D��]u��
��5o5��g�u�S�#��Ay ����!-~G!�
ς�i�����~�yH�%����sb�ɍ �n��=��E`i���p̉
�4f�؍�&���sH�4'�k!
����ѭ�����#2)�b�;�sB�EX��$u�VF�Y���J,�bK���v4n��t����j�O� W����0�t� %��]���s�եJŵ�o~����M,O��Z"��N¹�����4f4�#zj����r��凶��Y0�8{n�:z
Lfy�铅���i9�<�XKeB/�6�Z�7}C�<ti�mC��wOn̑��JZ+2��0���;p|I7�1��;蠹�rf;>�+r�	��m =|����kd�S@	���� �ڽ��BQ}&_�����Z�ybnLH�=x��ɣzW#���O;�5�����@t���ߜ\џ�RF� AeX{��<��Y���Pm��9��;i��N��b��"BZs�S���:����6�RP���~�A��`
���-��T�0\� ��6e]q�`c"�m�T��7Xw*�<r�Z�jLU�Р*3)1� ���6��t�&@G���Q)�b,=.�r����sv�8����xZ � 
�h�J,�:� NK��]~
n(0vN�	��I��ߴ���bQ��	N�'��-���ogV��s� ����R}jX9��uUM��B�#�v�E�U�!��eKq��;��(�p��n:��h,��	'g�MUP� �c-��x���X��N\{%Q�����x�B���R��ንa/h@q9����]���(�wȯz�Ę��Q �j� @���?�G�"�UWq�����J["�R4'��ʑ�PkZ��pJ��I�Rk��Z<��e5�w���w��|@�XN�"��	n�5�U@ɧ����@��RY�����.�����i$M�" ܞi>t/�����ww�J�ў�J�e��\�|��ޔ��ڸf�*�bDM��NM9��:oh_����i.*�<�`0X�#�YSIJ�o�������+�U䬈��L��P���QFɧ�w�D�����Wm� �R� ҩXLXt�bi�"AGE5 c�t��_�M���9���;ϕd�mƞ�i��?*0k~E��.���h��n�����E˹n� �����H&�BH�,��'�{���;ǉm�w��#0v�7�����io~�0}��3�|����U�1dXA23'���?dp�o�k��(BFe�;~�����\�[�t�w��r��;�)i�"��.�b8��~���/8`Vsӓ��U<c��#����#�m� �WK?d�1Q>&ԝ�1|���e�}a���ź�֯�+���0pY}��!��Ps�����,�1�*�םUQ����Л���WO�[��0��%B�"B��#5�������1bļB��7{�<dD�4��r�Hz��¸y�~.E���9L-d|К�lg;I�KF��J�h:��p�	<@-R��M6��ゥ^Ĥd�C�B����ϟƝ���*�6�$_ժ��}�&�Y�T%�2!G_���輖��n�N֥��R_�M�gz��Кz+����zi�kx���p�8�/R�+�N����X���j�T�&���򋯞�u�j�#��eof���1,���8�.��v�L-���3�W�qۖB(:,���r�T���\��B��2橎Ę<xaF��&�6 ��� 0:�'�����
�-��b��/�Y%�EO�ĲUBx���Z�7[|���*�n�}�F�Ɍ�`o�|��p�&,��ƗG�U�$���	I;��T*I��5�a�;Z��/�0��|󟼀�G�._�a�Ӓ`1�&jM;���Y�; 36�8�����Oo9��x�����P�Wr��W�0'�jDw���:ד����`��+���vh͇�RC��}���~&l�~�A/�u��G�0&��']�ޘ�� �]!�n-`�au�չ\���}�IF���� ���bLuջ�wsh��I�C?�M�z�2L��rՖ��ܖ�]dl�>aj%�Ǉ�m�2�S;&4a�&�X��W/��x�U�ߓ���!�@�V75	��|�Ar��V�>�%�:�K�hҎ91�x�=ᒋOkV��g�ԏ{\�]{ |�=>"�3��m��Ba&�`�oj��mM�dԟ�ħ��6N�̠����72��k&���왑~��
�Cx'У巨�,��׀��˿��Zs���;�$�H4�#��Q�j.$��c��c�(��Ur��(sL�t;���4F1yL�4~��_`�i�@u�{�N�kC��ܩow��Ն\��u6x.f��b`� �s>�N�֨{'�F5ZN��F�6tў`
�p� �"H@q1���u�{�9�_��!��;O��A�$� �����IK��GF�h=�m�w���5�r�!R3��Lܼ߸������^Dn���w$i��\R���y ��|6��"�N���U�|���	�x^U��G�$�?�L�mN��#��sC����M�;:� s�s��7/ϵ��xN4�����b^��Y9ٍx:�8�Ż����90-�]nN�y����SA�{�E�?܁��������0�}��߳����B���w�p�����6dLc����%ǖC�p�N%��.��^�W���X�!1�C�2��\���3'k@ξ�._S'q��c��c�7\�+*@�@�_J[���Ϙ�·D*wb�E��v0�\��6�m�,�a/��Yܩ���0v0���;{��_�Y���'#�eK���������:�p��Y��=cɵ��ToO?j,�<�@�M��8���q���I��������}OQgg��G�Q�kb������Z)���M{�j��� M�6̪��!$3�RW��]�G��N��6p��7�_�5��$_җ�(>���S�NI� pWM� �\�٤nȫN�X�e��ۊ�����qg�~�w�����~��'C��P���ON��Zv*�H�1�Dޞ�ey�e�]�qM���M5Nϊ���&|A����5��n���]�ҍ�����/4>-�#��}�E��D0;XGs�7��	�	��! ���t*�*(�,��$U@8����s��Y�!�L����4��tm�-�@\IA[�ER_�W��),?�3�ך�'זX0Ֆh.G��g��6I�o�%���'寊��$nY,{�"��=���[0�z���Af�fR	]��[cc)qP&�'��vR�c)T`NA���!�y �ٳ�������V�	 #�����Yg�oG@��f�E@�
Ʈ|���/�,�q���%���rp�>��ɒ�2_`�@,��}�齣��B5��	v&Σb ��ɑ�
sq��ؕ(q��������'��R���킑�>�A�r�o{�>�]��_�"��*�� �&
���V���8Yx"��
�oYC�UO��� Ou�A��&W,�#���^��!���f�7O>�:د)[���� �0I��O�Ӣ���lG����_j�n�=>ePXSZ�r�����ܨ������~���3��5�E,�1�܎dV[t0���ݵڃ���k�VH�%M�ڙ��m&yH5/xu-�r��#}�|�)�v�]�Jӂ�f~�r��g�i��V�m�</��D�([��O,%. ��]���+�����<𚁄�z=�f�:򣁥@5�&��]�GD����� b0�3��g�D���R������ik��r�f��!Q�sm+n��-K�	2�Sd|��z�.IЙ�uG�c6b�l%�y�`�����uVܿ٬�b����D�h�&Z�{����*��֗=�ʺ	{'��گ�3���h+|./��(g
� �+�0��(0}x��R�'�~�<toݵ��wM���1����SӶ�҇�a�qPƞ�j��d;��gЫ�*N9n㦑$��K"�_��ޕ�I����Y��� .z�j"���?�{�t���,:���4:�٘C�7� ٲ
x1�9�l�y�<��i��F��a�d��g.��"]�l��qw!;��%@pKKW���M�$迱��מ6X{��F���E����}r�jWLl�1�f���(�E��LH���ħ�O�O[[[�b�0s�E��J�w���{V#����������h8e�TrD�;n��¾�/��Mz�щ~C�
�Vz�L���*b��-�jD�!�}ҿ|����r���̋�	�TS�؆L����>XYe�o�h��@��˒����4-�C�v�F�v�$f���p�=�����0�AnM������ �r~��dð��W�K�
�Ҽ��RC,U��r#����HZ�OQg) ��K�xvi���w#�����?��ǿ���)��ŵˉ=�=KE�tZ�P�5�(F-���~�5a}2��B���@v���}����4;�9U��B���e��Aѯ� �O���NcO!a�����Єd���"���Β%j�T������}k&�~�z�9gN�(E}҃��~�ў|f�lzT|ڨA��1���%%t[�llU�L�"�6	�8�=��=���y򁏆�a_�Ά�`�/+wS��z��aӗߜ��X�L%͎2���]��YΗ:B����ZbM�)��4�da� `J��f�q�	'V�4�m˺N�E��d>��h�u�#P>��~2(���)X�/j�Nl�	ּ�;�s�9'����&dR GB� �Z��� *L��~��vXO���)gAV� ��.|w�]��S���J/��l
I���?�c��K��.��G5 H�$H��c���ŉ��R�&�	�8r�9�ܕB@��}�i��FǙ4�
�o��j�{m~1ܞ�7hm��6�������	�[d�2����A�i�сWL��Uo,o��rE5�0U=��cI�q)j�[w��R��9,h嫌���2��2��&9S:!�y&Y�?��|VjҊc��^:;�}e��W�\���E]��v�?|�$S�^q�0M��7�ijL��v2Nқ�(Q�<�T>a-���E���㿿J,@f�oaJM��*p+W"�"z�¡#���cô����I��ct>n�D������x��R�6#�|d�Ql��_Ƈ����臨}��	JdD�|H�?�Xg�F����B�O�{�j���y�U�������ϙ�}��C��H!���z�p�~6ڴ��l��uA��3���Au�R/�Z�m-#mf-��ˍuF�����'IE��M���rk�R�_ph��F��[��S*8G�ݸ�X݅O��9�"gE����]yk�4k��s��Ʌ]8ȃg-Y������V�&�֞���jY"�f��mA��T��?�Wl)mU��ST�X�(��V�l���7g��ҔS�(6�C-��4[����������w��:5��r�<����� �`jxv��@E�f�_$g# Rs ��M����> ǣ��H���hc|_����ly�0u{� b������4ه��Q ����ɉ�o�J�JB��/�?�|�(XKu��'(�~��b�^E�d�Bvz��� 
޺9}=�9��ok=���l��:h�R��}�6t��lԵ���L���Y6�JWX 
w�r�f�T���B�:���y�]�%���#��g�Q��}��f>�Z/ί�;���2O�c�E�E_�^Ϯ��~l���� �?��|�tAciUoI�x;quuZp04�����̰���u Oٍ	�,���@�@{�o&�����p�S�7;�|��2�=	g�4�7�Ϋ���|"VM��UvA?Y�f|�C>-~�i䂿z$&����Ƙ����,^A��2���Ć!�94�t޶";O�/!]m���y����L>�P���A�E����Nޞn��S	c`m���������(�ϯz��K�lT̽�T˃6|֗�#_�ƅ��KCwX��Ew��Dd�͈��y�)�N��N��j�����Q.eٰ�F������`����JE��*Ž�N
Ei59�Ɠ�<,��i�^�}��z�r�|���-�r���o�'S1�'�I�×L��Љ-�~����|P���7I���i���
_�"�D?g�e����q��ߟ�>�*��dˊ=��L�
t�n����]ٺ;v�y���R�ǥUxp���r��3�R���`B��`�zĽ��)����6!{}4?-P"(Zp��n@K��7}?NI���J��\�>�C��Z^�# �7F@b6�4R}�^9�h�j�O� / �G\5�qu�?ʥb��|i!b�དྷ��;�������'���؃�K3��mU���y��#Z���]���Ӡ�S?�}�;<Η��B���b�#OM���Y�X���Hn���"��''�����4]��[��1�ڛ~����E>�7�P����ǦEN�Dįb�z9~'׬k�{��-���+�	y��_YLջ�����`~����º�o��V|���T��;��"�ـU�l[����=���,��	Hh���!80�BR������3��u	Էv]�~��rU}/��y^|��&I!�oL��/�m�h{�3�#H��0f|s�̘���hO&��lh�'h��&O� ��I�l4:`���8����-���4��f^��S��0�P������x���@λӋ������&i�E�I�UG�)f�М�_f��$�T��_ډ�r(X����1�1ڵ��1�΢��>�_t}�-"�)A64���e�P�C��nq�M�0lu6	��P�̰	I=��J�Ā�ěv��<B�����Q���w݋��`�b��F�'t96�^+ߑ�WJz���!� %�]?���j|-���R@Km�J�F�Y�x�`��C�.͠"D8�J�ۻb��6Tǅ�� 1�����4;U�l�+&h���x'�7���2A��q�_�OD]�B��&��a:Ƈ/v��¢��~˲v/�+7'k���w��n}�E7W٪X7s� �E�Φ58`}P��dʽ�jT5=x��` \�MR��IJW�2�U�7B.�|��[��0I�ϱ�F1��4�4ft ������G��A�Z#���-̿��D_����ƋuLVl�Ю�]�n	�������>\�ח S(s邇:ϵ^U)�8�������9�ֿͧ�M��:%��4i��f6#a�:QJ�j�ƃ�j��bD�Z�c��&p!'mz�X��i:"��� �3MdC�F�	�O��;�\���x66Dh|ڥ @�Ae��ī���bm�|IJ����W�%8�?`@g�42��]� '{它� �=���qƊ��Kؘ`���	�	9[��Q8�Ҍ�ly��W{;O)���|x���<�]Ϗ��ń����*	I�!�������j��Z�E�ٍZ���E������퐤��ܹ'Y���� ��ơ;?��z�V�{�Ů|���A�;U�~(<},��ٞ�b�utYf\�:s�~��M��1�
��PoX|)���9���D�##&�^U%=_�ڳ�?����q�%� �9�%A��7��,ݍz�fYɺg�W�q*%|ԩ<`����<'�<B �=�w���*�`Χ��T��I�[�ϝ.��?yq5F?xM��9$��p�Ρ�zT���U����f}f?�!���͸��Vw��L6�z�_|�N���}��ᣣ�.�o3�AmT�^7K��R�#�X#Ώ6ogO�\o}	�2ïl��(>��r�B;�!�4�ND�6M�gc�Z���y0A^��kF*����md��!�F��;e�/&��2ks�LJ�i�g�*e���,֨�<�:Z�� b���ű���=�Դ����U�zLL�83�ծ�QB+���ab��x�]��|���?�/���V���`ߛģ��rudvv}��0U�Jf�I%uH�Ք�h�D�(����iR�lY4�l�Y��A�5+���P��7��rꚵ_%���ź�KӍ^"���h9O���>���1���)��D�� �:�����5�NHxWT�p"��(�y2���޵r+���}��o��*��*pͳX	�b�rd��]#p�29�������$�����܌��/K��!Wj�W�I�V�?�tz��˂	\/Jg�K��ܷͿλ���l��ވd�RV!�x�����/�(cF�F��FV��J{ߨT����:���>w��щe�G2svG%�!�
���"2@͋\3�)PSq2@T�I!���6����"�دD�1�"Ya��� ���+,����`
(ٕA�P{�y�izwyOE�������+]&��y��+o�"�1R=����=��#���1��i�z�x�B2A���x�=��^�6u8�g��<�ZWo8�K4T�:�3:��,o.bE��-~���Æ����m{l$�1�!㛒��?���ă8��fD�}]�To�4A��ݧþ�~��|wP&
�����<#AZ#խ%cM��j��>�F,
}�+��]xI���; �̈́E�~u*��&� �9z�u_܊��'$����G"�X���ɂ밧�X��B����	�4���i���F��v�@Ӆ�8p-:�xq�~�[d�X|+�b��|�2�s+�6-��%�iB�|�{�"Ǳp�Z�)��S��@{���NHۅ�`hT���QaKd�3����.aҎ*.Q����8M�2}�U$1������9��v+�#�7C2�L*�:"1�/S�B cm-*f:�v�)F0%��j�#��������R��UTZ}��v�uӽǵ��A�}�a<�x���Z��gXl���g��x�EZ���vW�I�	#�ҙ�Zw}�LB���������>��]��K����;i�1쩣�Ґ�!�"M��s�(L¡����3Q!�_Q�	�"��k� ���Ӽ:�mx���l�}Q������zv��W����Y�dy_�鳕����4�%�3hoE�<����!���9w��D��\@���}-�й0,���+s�E�:����<�`���c�[�4�mZ/���gT�;��\%��O�gr���x�e�>Ɲ&��=X���|3��|�t	�/��v�#��ޣV�~�]�=|��bͥ�qv��=6H���s���m~�(0���-�k̝���`I��-�Gɏ :��{<Uc�Gk0���r,��!�b�g����[���M`�x�b�Y��^�b]k�ٍh�/�a���f����B�O�[�mD|x$pfM�7�폿���Ǝ�D�9��@��(���%fN�j�IX�"K3|*���G�l~z��p�1����V��@voPe=a�u$[��/��䭶t��܋�hV HR����
�*u�>��bQ[�`?m��쒇C��x�qXޠ�q"H�Tu��!�y��&�V3�D����I�����Á�?d7�8�,8<v2���4ފ���D�F�S� ֿ� h�ٯ��*�d~�R��4c{�w��'��vӤ	�Ȼ���86������J�a���O6m���3%��]�C3e��n�L�qZ`b�T�[B럥z�Y�<>p�uWM�����XW'7	��4�|�w	�r ���bs�l�?99���+�SS��<�e|H���=yܳ:�ߢ�Ew�qh����T����H���Сi��_ƭ�·p��l�O�����Z�{�U_�t���15�F#]�H��J��FD �ҡ�0R@b�t+HH#�"����y�����v8�����뺯�N���J�i�BJ�G�"��&�y���]-ʈ�%D0�������:�w��$~�Q7x���hV9!��[�p`ãC�I��0�_�9����c�炙\��9�P�I��a�����(��0lrq��\a�듻�
4��mo0���3+ L������������1�Y�"��]�}q�X�h���T����}�.�B���Y.�<J�E�Θg�����Q����`T��
��ӽ	/ԫ����h�g�H�c}=��l�H����ޔ�ˇ8p�
2�����g.��Z| j��_B�Q�H՚E��w1P}	��D�H�}��6�-�f�`���oև� �t�d��s.p���!�}ϋ��S��Q'.���������ڋ��rJ����J�p3��
?�E�GO>���� ��{����t(��CI� �y�V��å��k���6�kk��>R��֨_{�?�]"B�L�#�9�;�<;2k�N�N�beJ&�ww��@>�4z�$��[U�+�*���a�y�ps8��M�r>�Vad���F�f��{����UDY���)I�#&}5w���E_�$�8L�s9"E5y3f<n�&G���o����~F[=�c|�9�ա�@�XR�'�<5D	*��F�:>��Y{?��rǀ�ϱ"�I��BP0�u�6�?�������7ֲ�������Pr��L�u0U|c���_�ޞΘ�����x�c'ϳ=��xH_�a F���p��wd�ꁜ��t���U��Ƈ�+��VG'\���05��-)ӯ/%�"Ud,Z	ﶄ��l0-z�.ĀE�d�p�&����&��?�0;���=~��>�9�n#i��eÿ����$�4jU�?K��BU�^£�_�i�A�S�!VWA5L�y�5�JM��,]�'o�4
��=�L���\���a��3�s��W��*bIBj�&y�S�]��\�.���(�;�3V=ٲ썢�:��	}a�9��юḿ��%��7c���Bn',���B_��٣J�kN��~"8���ɇϋ�.��H���A �O6���c"xD�1��ֱ��0�zMZ����3m��Eؚ��ґ"̃p�L�e�ZK��/M�x��s��r#V�EbS�Y��_�ӡZ��A-���;��"�P�"����L켝�;3�j�3�;�!�2��uv$��|r3ߔ�K�IV�X�R4�5&P�����n{}:JH���9�^9`rF��k�� ��/�"V�=	��/�,��|��������{��+v�;)I��X�{��8����2�ങbf����������#�����)�]f��<� B�=V>��=qRa���3��
��V'V��h�t���DpWs	J�* ZL����]�q�0��݂a"^?�p��:���V{��MFrdf���1q��:��4���B�З-��ֈp�<�$��r�uv��W�}��4oAD��� �?�L^n�@�é�2 7@>!��#Bw��� h^B\���Awf���5P7͟����B�+��
q9��9>	������̵�U�e	6����ck�ƕ�Gw)��M.gN�F��.Bx Nak���M��,��@���#y/�k.1D����z�nbD:�֯o� >�4Ɍ��F*F��K��!��-g��\��>r�7�	�j<��43�_Cw�t�!��٤!��@�p*��+��KR�e�l�w�J� �y����?	�나����.!���b�������I�f��]�� �;;�4	���r>��%�J�{�J�o����p���x
4q���y�z�0�CvU���~y�'I����$Vw#P��� ��V�V�TJ�q-���Pj�#x����ԇx��{3�wS�X��(,��i"�>��M|k��ſt�&� �0i���{z `m�&� %���f1<��ic��rE�����Ι'G����Y���� K#H���GS���\�=���܆�<�#h��IF�N�iFaQo�s!���)ie������g]Ag¼��Ӯ³�+��:��p��a�oI4b�	�s��^E��x"���a�t�HW,F�^�#������4au��|;�U���(�֝�����\��3[o��訟c���MW�J�m2Q�Dh�6��!����[+n���] �?�q�k��SzǄ T(,:�Ԥ���`�;�d#{�C�QWm>~KHo@��i�hP���BD���Y�:����B���D:�&a|��qf�w!�������f"Zi��07��<^{L�|�������& �Q�+p���sP��ԕ��x��~|��a�����A�ϲ�x�Opa�ƺMV�F=�8��ӝ���7���z�-.��܊Cag�������+R��L���΂w�B�3��l5�ժ�I�"-<��]��~�5�p�v{���@��à�[��V�?��X��P�S"P����0܌Q����y*�ޜ��s�jI�dbH�%����do���:�e���H����3f��$� �.��?H�ve$N�~��/N�	�wV�_v�OV)0������vQ�����吮v����|�'ݪ��WV�`*�MƪR���z;���� >�_��)h�Z����g���4Yy����5rek��{�
)ԓz���؅$�����ܑ�R��,"*�ԡ�H��.���{�b�-�t�{ҍ�B��v
�Hn	5���\�C����� ���+�{?').|b/�\p?Y�E�8E51����0�ٽ�Ţ�Q���1�R���kp���.]Vw������ߑw�'�q�[�ڄ�I��;[߾�{�	�¶R_�
.��_���xL~�}"���1���,��Ҙ�j� Bs�����W��D����-o��$������zLf��}q��eH|��
4*����&��4q8�#P��<N�=�'�k�p��5,/�٥�1=��awI�2�H�^{gH �{�{�P�>���i�X�X�ݻl�)s���$�f�5��g�?E*R����b�lU�t��CD��z�R�����c��	&�{Y�~PȖ�Ì|����W(��ؤ`fPg��U�>+c�1A!Kʮ5;cb\oC� cʛ�^"Jܷ*}��@h��B<D��&�@ ��������)J����.1��;�?\`y��£e�[��U��c!��Y]O�67��\|O�#^P���'�p�ps&�#�T�(ǲ�v� s��Q�nQu�t��*��� V��X1�_���N��U�zM�~���f/i1��Kz�s��˨x�A��Uz���WQ�,3���F��,�욹�I-�Y���W8uj���Zv�\��4I�ߢ�E|��M��#W����Wm����c���z�$�Z�H�³Qu��_�B�j�`����ߝ��k��2�����+�� xVZ����H��*0W=�n�Z�G��Z�b}Q�?d�@4�qJ�CFD�Y�(>�r��D_w�'�_b:e�62׽#ch��W�"�J�J��ޡ6E[��'��|�W����ן "s�m�z���q�M#���3f9�����471n�����p��A��$���g�dH �WGo�]�)$FRD�v�v.A쎢���	~V��B��`f�e���m�,޹�&�с��k�~Zym�ʵ{n����^�Mb	�������̛5���g��
��N�0\���0�~|�'K�XV���(PfБ����[���ʅK]�}8�/�T�a���p�������)ez�1�Fo��f&}��������P �T�M�'���^��|r�?�������X�����t����0$x��==�Wd)�����Е�W�'��|���!$��]��҄u�&�<Fr���6�!b��%6dur�o,�AJLD��H�#?:U���L���3ˇ��*$�����"��}Rsۊz3R�Vl�UD_.�+���?��!L@���Yt��e~���#�ȏ��c���rz����»jSӌxĂ��+��=sη��{�hy�7��ڜ2O�+�ףYu�{�����g����h�U߇��On��M�lOn�	���_��L��Ng��+tu&VS���Sn����H(IƂ�Z3�����UG|u5�ϒ����Ĕ��#�����\�qX.��������g���޴�~u|n»`��13�֫A�}0�x�D{[�a��t�f��)p�!��n�>�q`���߆O�#k/R�̤@� Gk\�>���j��ޑ�U�-,�KI��Z}�~��d$K\G,�]6��yh�hQ�:9I����y�ye��g�����p�%qԑ��<�� B��fd>F_Y�^`�38G�!����*���¼Y��m'��xOI{{]C�魔��/Ї�uE���6��Ec%��
�=�i�	��heN�}� «�RΓ��n���!#�I��+_�B#����>���Ի���nx,�oV0�i����*�<�d7/���K*������n�-o:�ωߊ�-7���Ȓx>��^̑��$
k:qG��(҉�gӞ��ڬ���MϘ���{o��y.�<�F���Uh���C����כ��Cf�d���<��I5�x&��>�"�A��������I��։޴O�&�#ٕ���{1~yAJ,����^�%���$��pD�@���ơ�m�fz���jO����$���굲E�~�QEb��"��;���N2���*�~�קg�k:G	�	� ���۸�E����h����䍢x���e����=&��QJ��o�k[P �.v�C�ήR�(�X��J��X��x��#�p�#hܚ3��" �V���*T ��$7�@?�j���Y����p�ݴ�}0�u��aD�>����I�ˁ�^Au��SRD�-�!e�e��~ǵ3�\a���_������}ɶ����*|$��6��_�2Kn���q�/�ٝ�[`��dZ�e�D���|��N��7H�3+e۹�����t�#�r�xm��<��Ly3��BϾ�J�w�Ρ�ɋ;���ύUp��Τ>��--\����b���3	icF��I�Rx�4;Efٽ�ĒX�xL�s^�u:�z�R���-(P���y�*�؄�0bN�-,��=�N��ձ���Çl�8�=p���S���_�ڍx�����dKޛot���t�$V�\C��),3�Rb\_{U%�`0�r�5y߸�'�4k	z��p�n��@�h͋H`p�G��zoq�7�Sdo#���c�MJ7Z`v�T���z����C��ϗ�L[8�+��ȼLw��P{�^\�)��c~1"wC�^��G��g�=��IHϣ|��&x �{�igLϬ�Ov�j��B���Ɏ���)1��F�_��<���,������S:���0H�X-V����һK�eרβ=�!����a4�q��27��?�r:��yA�Q��0z��o2�����𾯵��C]{K����3�ʟ��
n��g��ç��?2�Ii�s��l�#�eKe�Zk�_�劽�M2�\]J�1�I��o�(��4��g,�;�߼���$��.�턨��Y�Od�Q�wm��0Ȏ߂�S�2�L�� �w�g�Š��u�,J\���ѻl�]�$���:�<���'�=�|/gi6ƴ�P��n:��^��������M~��HsV>�~�+�J�K�^�Sv���[�D�y�H�]��"�*'�ҵ�J(����`?�W�Z��e ����r�Q�~U���q�n��|M���r��X�X��=��t�|�X4�3��b�&{%A�>�V�h;�nP54f78/�"�F Ê{mЬH���v<3#��Is�6���z����ќ'�1L?�a�$CקFh�;%[�cȳ����a|��ꛬV�p�� �[���Å���|C�쥎�������:�vˑ�����������6�c�lcQ�l}Ep�⓿a/o��LO��i���
����J��KOZh��]=�r���`=���w���Uɠ~���S��C�:��W��u,�X�N"'�u)N���u8޼� ��WMV;�E�?���G�5�+a���Y�4#�|��zW�!�xl���o��6�M1&]�㳏�S���zw-��? ����/?N���
��$�HC�$��1b*U!��)D�  (d��4Ig���{�t�^=�bL($J��w���r��L��и���T�_!)��Ê��Xp`���h>ݡk�?����2;�e���u����pY}�xY�]��@�fɣd���S�`oHp�JP�	d.���nfpEc�3����EI�(������8�)�[�����Z����:����恦�{����ϵ]�H.z�puH(h�@B���"�D=�~������ӯr�Pqm����I��C<�rFj�;�~o�#�|mF_];V�sR�i��픳?�3���cc$NIz�����M���\������Mj������3C&3s͹��v,��jd�Jj����L��5>�5��=u��^?/1�rR�\l���[�4|>�
2j��̓{=�}��!W� 	X<�>J_�e�Ηs����>h����7詻^A�������M�<�~�>��Y�WX�jڠ#xr�צ�q�g�(V�IE,�'�d�D�� �3^(_,ޯ
������c�og��!c�Ċ��b=��0?齗�+SF�YZ�L}��������K-\�o��"�n�c�MYtN��+�D�g�ZM�����F��uŸK�3�� �Y�N>!=���6���0��� G�<_K�ʯ7,v�ߞ��ܞ���oFzn�l���Ls�9�`H	�d����-�����N�ſ���l�� lq|�^hӶ5B�
ˏ�?7k���e�O�b��i?��S�\�\9}X��3؍��Dl^� ax���yj��	=鼱Ӣ��\U������vO�6���6��ѫU}+6�Hү4!^c��� ��'�'F'�\q����\�uO��M���%6����#&�V_~K/g���d^�^�H�u���״�;1^��;O��=�E����M0�����þ\�B����V�=��T:!������qM|'zTD"+��HиAS�|t��ͨw�6xN?�[�+�'�ߞ�f����B8�'���O.�]�(�_Ѿ�E����z�ʼ�����/�o�PD�L{��?A���YEeAfH���GDޚK�%�p��bgF���ɴ��3$7��o�EV>����m<������
��� ��i8}`��|2D��ip>!�Y"s�+cbFG���a_��?4��.�<��>�7����d���g�|����W�4%I����Y��pA�Ⱥ���#7F^7f^����h�[���}փ/���3�?]0�r���szu39����k���|,���U��A޷��L���m��5��2	��W��݉R4�k@�/+H%2�[��ۀ@?�zT��]X3�E������T5�LH�"���} �� �G��!�f��b�US��&�v��G~jeK4�4'}��h�
�h0?�f�+�sMA���&���qF�Ʒ���D>��j��;�� 0�R��δ4��%��XY�,T�% �~ɇ��#Q+��h�E�����>N�|�1��8,	6�6Y&�5\��.�K�Zr�mQ�0��{W�p�EFZ\Q��3�i�:$|@��/�(����V��2�6�㦥*_9|��DgH��R�c���6�m2�;��?7��lFj��3}P1�W-)Z����f�<�Z�3�-���r����y~]�
+�N��H�/~�������\�����������������vS}�lͲ���ŶXm��^LP�G�n��$V_�]��'���l����3z��H�*i�:�k�g��>�`	HgXH��}�PF�z[j��kE�Ũ|��ސ�
�*ԓ�o��7��e	�j����_]h���N@��,�-m��h���Rڹ���!J(S�cVp�ʧkw����C�ٻ��R������#EZ=�B7oc��G�&	H1���ϨΌLɿ��E�#J&� |�qyMTO��J螽�.Ҕ/裱z"^	G��x�C~����Ƈê�H ���?�yD�OΟ���^V�R20��0���_�N��^��y��X�x��>�<��Jcv9w���d���V���Ճ�LV��{�����ѾiAi��8�xy��P'�
j���wF���YYv���,����s��y�-�/]"�.M,�Ç�'׿4�U���pX����UrM7��yG�u��o���E�oH~���J`�y)�����0?I&��m�.��Dr;�q�l���F� �����I���;����MX�[�P!�niaDdm�"��@diuNڂY�	�2��15���O���a�p��%��]?K�t�O�:�	A0�\�U~��n5j��7Lq���1@�&��Q�J��W �v��I�H�.4�찴d4�W�E���C���	_Nq�	ubQ��{�f%V���O9���Ap�Վ��Ym!�s���w+(0z~S��U�bxc ��dl��F)�ה� �o���������P'5mL'-�N����*m)���H�����/k��m��cm�L��� ���5���$�	���"����,c�z������ZՃ��7�k����/&��D�>)ڪ��'.���� G���&ك�Y�zFlT��d����b��^���ue� Q�����hlٛ
�~0a���l�׾Ď��	��ާ2� I�|��"G�{�[_�<������M@!ؿ��,����y��:p�$ �#�Ai����@d��.l��G�2�9�4s�S���=��.�^����8��Y|�YV8t#���ݱ�I���n����/Gm�
��sr�L�4,W��Ѭa�$y�ylP�䪉ִW����a�vЙ_�SR2���\C�����ʣ+}�����J��
��6�+�����֊���"��,��Q���ay#��c?��S��e����z�<����Ut�=����Z�lM)z��nDlY|�����A�b���CC����z����o3_�ˊ����i���d����CAc�<B�PZ" ��,N��������-��u���/��Є��k��n��*�U�=��/a��44�\�ܓ��#�DX2B�{O7�K�T~�j}U&�x5��Mf�7�J����1޼�q`�<H�G�t��K��F;����C ��ƌ��E���DH�A!yi�3����2,��aˉ������yhw���I�8:�q'��u��"����#��K��u��=�>c���_C��`�Tht��W奡70��jF�Z�#�?S;@�)Ы�	�0YB!��Q���I��s��}�'�?sF��Y.G�|�כDV����L2�n����?������n��4��e��]oG&�QC�����<ۊ�[V��B86��le�MZ8�|r�sN�<�ү��I�xW��� ٿ�ge�r�+Q)俥����ւYE�.#AD���P��x��uT]�E�9 j�w8s�;�:�w+�[`4� �m�����:?�S"0p�w�d������D,d��or�DSǇ�}v͸��ƞ5����Hΐ���?+A�L�B����n9"�q�����~�)Ȁ�xXW�<���0gQ�ȘyR�oZ�ا��ȃ��t�0���[J��f8sT��+��Pɳi*�݋X\�Z����س3�v�U���I.��!�Bc�g�H�	P���7go�\^E�挰m]e�K[�[֏!��w=~�Z���N�����	ئ��	X�����}����YG�2�	��0)���?�H:�X���G�Z��R~��mc��*,��^�e�}����Bsx������XN �2�����t�1�y�uÓ�xR��D��{�8W{"� \bI� �OF:qR��`c#V̥S	<����O��og�F�Q�~e�^�wײ�q� �l�n������:U��µ��{�҂u�t3}�)ͪ���� �z��H/'��d6��sH�Wuc%5����m����r�O��Ѧ(6U����uNw{��߂8A�^/�������U��8�{�@�@�6y"%jO83�w�˭��!$s�o�ȏe�Ph%>>V����>�$��:����}�hJb�����ϔ��0�_OiD�ki7�w��f_I}�����r���z���"�c�0O�e�a���u�£�c�ۆ�I��AN��8���u�:n����g��gpuZ���V���#�9�{��4ٖ����MA���͙���\t6j?�Ed ��o��~n0��0e;e�C7�ѫ�3�bG��|�;��m�����!���HP�и2�N�6�M}߳Pֳ�6���|�64u\$�b�DB�v\�$=�*�����q�57Q)��bƈ��"��l9��jsA�(5�����Ĕ�&;oXU���G5����'���]��@��Y���'�M���� �G�0%�f1��pV
��#E� �o��-#��A
���3��H{*E���!�}��Պe�}��w��}�� >Au&�ze��2z�X�T͙�x��m*,}�e9�RM��6}��K}����6K�}����m��wy��:v��l{�-?���/2����� nL�seỽe5L�O�D{pE䯩l�p��L:[:(o�����nM�����(柳:#{��&H�m�����5� I!H�g�ѽ��(�Z��}0�B�7��\m���F��;N��e��u<�9B\��:��%�1��C7gЗ�.�^YaɬQ�\���9{C9���pD"G:����&e!X;~R�<2˹�;1A��\N�~�4����B����MS�]�*�>/x�(�kx�}/i�}5������p�����]KhEĴ��m��L����-����6�1_�?S�r���S����Z�
2�o�M��@��qW�ú��(Q��8&�9۰���v��]���w���.�mR~O;"���M�]�wױ��3)ޚ�KSF����4���1~�������J^S�N�������gy�b?���L� ����L�2Ok1�n�J)O�����cE���"I�rԶ�������,����G?��ٗ�#��"�w\����Ŋ�S*&�[����8�e�����5,i���WÞH3h�ꂆ#l�	���!����M�X�|+R�y�o�~��@%�ގ�!�@e��l<�C��'��Hp���--���\�cHR���ؗ���+8i̘�~;6z���Do��3:���f*8F-�����4�v�ަ�L��|x_���y.��뽚=qu������0���Y�	ێ�k߆��� �έ�	|�}�S�}U�[1��،}	Y���g7��X��柇�����]8+>y(/��勿��P�v�ظy!^��ܴ]�|l��O,��ۡz��O�_��#Ȏ��[$z�ȇő[$b1�����]���^�-�2���0�Seo�<0��F@�!����n���qn�U_�Ԧ�6�Sk�=wszQj ˌR-���ˏO:ĔX�g���= ��@$��Y&J,�Q��5�d�� �J�J��f���A�N��7*�q�+n����9��ߨ��nYY�)]�?�O��$Z�<����6�*" ��Z���H������lz�d����J�wě�~��akϦI�����y�$�̣^��e&�]&����K�s��LEM'��*6f=�qI��&�E_]�л���t2QK��?l�(���џ<�UoT/�+�����ԕ}�D�Ev��w�T�3'�$D���Y�T���˾�C�% ��� h�YT:9��[>�4�(��Ue��ʥ��~bsM�Tı�Y�.G��s�F}����a�B�������p+"�8�	>Vc�t� j����ν�(��g�\�%���HI������F [!���=���(�[=θF	X��d������!+i��_��j��Җ��0w�W��Ugp�Kc^d����
�h��駴d��H�O=4=}�3�\���za_���?��]���Ec�ڷ����a�|ww����q��b)Q�s�7�����;&��%�'�z^�J9�2'  ��X���뢱����?��4?%�����+K�jt�|ҷ�¢����)3�l�`�#��nQ;dKM���`�F/�3k���*k�`�,�hj�*ח�3_�#�I�����UwӔ��ڲ��`�g7�,U9���}��>a�6zK��w�Y7<;|\&�7�ʶ��)��-K$b��JToA�����Tٛ����Ys���̈B��=���~ {���^YCjX� ���Z��"���`V�i�q8Lک&��qn��T�[T� �>qP�-z�>妊r<��G6��6�7{�M���y~2p6P#��D ��<��_�f��nE`/M�7�B�����Uz��|)��5�ԙ���2Bu�qjN[�F��iN���W�x����ߵ�_{�-9a��n@^1$�4&]�PM����/������C�Z�����+�F� ��o�'����D/8���l��0J����`~�ӛ/���N�����U�QV�O�~����Vvl�������R!�O���5�m������!18+Sm���9o2�f��n�:�:b��e�����Nvс��n�4��l� ��s���	���|v��&�W�!6n�1W��Os0Ŋ�d���3O1�& gۘ�W<Q�P������i!(�HNıQ�ZFըX$a�#��.-ʇNH����K�
�Ԍ$���~�W�0���9=@7��x&��Q�T�>Jgk(L^�mM��;�DD}yԽbjd�=gr(�:_��&n�b�P�,㤥����T����'�P`}*�q0�<8�?�c���IV���?���:�~�/
8U/L`P�P�,s�M�z��
ȟF�.&3�����6'���)�19��2�9O��B���/? q@˸�z���+2�1�z�̗�l��wm�Ң�P���q�03
�k#��D��O]��p�Q�xI����)n�C�Ήh*��ȥ��J�}UM�;C�Y�{+��!bza-���0��h�*�kGS��79,Ä�b��y��j�X���ω�3n��j@�b��zL�G�?4ƒiK���C���-`��꼱��D���NV�w�a�[��� ��=V����D��%Z��*�ٚo�o������X1{p���K>�w�Z��=$VXt���/������#;(\�]��|Z{��<�&b�um1�`)�SD�`s�Y�K7y�SX��EtxHpÎf��w���Fn�\]�̾�h�9#F���u��)�K)	ʫ�����\=�J#8� )~���r�C��O	D���G4��:�Ÿ��2/�����N� �Y��Yq]���0���
�&%ڎ �!`둴�0'�nzp�����*�2��𣇅��齼[Q���jCX�L-�C�猞�j(Q��j@�I�4��;��Co�C�8������4G��&#H�U����gC��*<��ǚ�����T��^���V9��l� �`:�|�ې]�]�ݏ�X)�Y��h��m�UQ�fp�)���J{Jڳ������A ]�E]Tޝ���v&+`�F�oXԊ\�_�c�o_� �X�������-�O�
�|oq�}C�kɽ6=*�l����I�n�}����t�2���_vx4�T',I6�|d���y�$��9�3�F�wL��$!�O������G�~KPÓ`FO6�_1�/����)�x_�P*{�B:�3i��r�H�&��%ʂaM�q}�(ˏ���������8�\[���`~0H����l��zm�h�>�3c��/���3~�K�C��m��-Y5{��������8�!`��|�6�{hͲ�p��W�eβ�n޻�/�o��J�j�=�n�p�;1��c���~�	��o�7N�ʀ��A��~�8S���F�$oK���ϣXb��9�[ף�/�}�����穋U?Ǽ�Z:g[��!�W'�҈t��b=��E��Gg���B�afB�K����N8�����K�6�_��ʟj�?�����j/y���o�Y�r��2�%�t�'%$ju������e!cTjV�����[��0��#⼔�Q��ku��bJӯ<�}�_5n6%(H�U����S��kpU�T��Z�J[�J*Tx�
I����B5�>l2c�K�qt���@I3~L�)=���Flm"����)6qW����DB '���+�E0�U�����63�g~7�q,��)������,w9k=A�+�X3�ճ���H�C	Q jZ�����Xa`fNxy�8�w����x���bdk��~��i�&~\��ћ��*�Y��g�4ڏ�s��#��g9p�T�&�t|����%yI�ܔuI ��ߜ��a��/j#�d��R&Z���f�V���N�!�xR���ef�N"Vƫr�!��A�}��*d�����}~�㩏s�٠W���~�����B�u�C7@�m�3O ��L�L#�`�FJ`}\��A���2��� ���zv4C"�}��mq�C|�	��2\��_�EK��rZ����`��� ��jAR>(0�H�dL{�/b?�o��F��ٳ�-��w���x�`���K�����_º���:��V+�F�XF;��i�����Q�E�p��������D�ߦE��8�
c�M�C���w�[�>
%	l����ڜN1?o��l�ڗRe�WR��^������9�_*�s��ޱ��z�G:�X��
��_��˚��|�d��Yx�>+��+jh�-J�ӚJ�agҤ�#������v�}+_{�Ï�����#�٫�����A_#�1�2�Ai!�$�+��9[�Rx�d���^�T#CC���;��nUt��2�����Z�G�0P��ʙx�Ąf6�1#,��B2�n(�f�i��lc�����	��~���l���&;h�*�`��,9�
�������v�!!bJ�  ��.#sRL	�l�g�\��O������(�^�&�`U���57Q��fz���4͡���z1���sFe&�Ⱥk��Z[�ݪ	8d���! EO������j�:aǬ��v�y]~�}p��5m)ۍ��J�k4f�(I����n�֑��պ�i>�I�?�r4v��X�f�œS)>��}��P�
���қ�4����t1���G�[|�_x���[ܽ(r0���`�|n�C����ˏ�����L��._v����G�!�V�(I\� �`X9�iZ��ሄ���n��F�r� >0�+�\'Gz#�C�<�n�[~k�{��SR������SMY����wo0Ak0�`Q@�,�Y�T�I����o�]7�*n��v7��`a-���w/�b���o|�_����k��
�87�S�8Qɘ����5=���'=�;�/�T#�Y��#��S/��RB 4,��ۑ��-�8��b����%

����hn��H�ΐ��斴Mѱ�5?u��q��TѮۍ��3�쁩��]�ğC���ݺ�3���&�L��P-�o�'$�67��6��j��gΎ>��9?wWy�OU~�婋K�?5<FAd+���.컭����������T��SS��𩫯����ro��1:�XD-�]�=���8b�(���I�����<U6�� 2ig}����c��f;�z7��w��A�=X�̛�m1�}��E�Cm���5��v�2W?�F;Ţ�xz�Q��긵������nX�،8/�F���(-��`���"M��5��>�q4��\@AB*ߗo�\�_��Ew���6��]�k�'�:D=��C�%�A7�`��`|O���7�H>ӽ�="I�Jy�!*�?!�����c���~, 76vU8p��5�I ���w���Ȅa������4�Oq2�}�Iq�J�%H��y��P��~�����eG0�g=��p c��˫�f���ӧyd�p����Ɣ(���v08�5�������Do��S�a��tM��ǹA��o+���o�2CC���5._���m����~��OI~�[�^�>��i��czE�'�	$$���oۙ���c�4��=�^�i,Tv�H'�S��?)I���ԜyƘ��g��ps&�k	�Y�c���	��t*��n�ɓ�PS��$t6�~���liF{a�㝽���G��Y�b� ͪK�Y�o ���ak��I��S��m�-�L�+����P,���_<Je��=:}���0C�e%��ٮ��1�y��m� �	a~KBSJ�gZ�h�Q㟹��#
�\1���,�� �[�>��WQ��,��������UC�<ܐ8kL��(m$���ۆ�@����+��NB�c��pKX� 7D�ͧ%!F�./kl�>���m�=/�X���+|�ԔL�)��g��+ׯ���c�o��*ic�9h���2����}_=ж�ǂ���@G�X�
�S��9[�i[��޲j0%�mR˚����@)�KV@�h�������G�WGE��_�0t7HwI� �!��)��9� �� -)-��1��t�tH~ý��~k͚�gN<����w������=v8!J���P��,���u��Kv��˔4eR;~Ϥ8�:d�=���+�U�h��<�D 1���V ���Rl��S��7+aD��x�u�NC�h�g��{m��q� l�c3�)�C[ep��H�?E��Y=�k�S/EP��l�A1d!�k���=j�8�n�	Ω`�IAe�W��^��.$161�G���:ëw��w�HIc*�e����l�~��a�YwԸ_���� w���3��(���ё$�des���P
g2 �,�v	��R�3�6�^!LBC�d��n`aЂ��0f房6Tx��@���glJ<P^I!�Jyd�4%E�uD�|\�p|��ln�p�"f��g���e�fJ�b��h�6�냮�f����9����K�7���e �K�d_���@~��	�6,Ncܬ&\�J���P�+���V��pRt�8�������e<������ֱk��B#��.%%G� E5���삹�wP��N�FX c�`N����_!�̴�Z��d+�ɵ��O�/j͵e��78I���_;���� �gW��s�����wܬ [���6"hH@W"�&��LT2-��
��RB'i��.R�'=�,��+ j�u�����ii,U��$��N�������jk�P�q������N������c����|mqb�c~����63]Nr���(� �U6��c�!2{j��aZ�!a��%�U��pY���޸���0%��*eE5��1vJ"��)Ղ���2ָ�J�#������ͼ���~�[�+Ų�1(��`�2e��m�pS�d�5���^E�}�E:�|if�)Eu>}
 ��\�}[n�Zܥ�|z8j�h�N>���� ����E[����h҄1�J*�
Q����}k�o�b ���%9�z�	���.:�a ��IO�s��H������&K������i�/Q�R-Q�{Gi�3^5��Q��cR��~�����^d�m~����N�#�?M3����'�g	�㻒|�u 1|?�6��d���x��N�v���e>��N�wR
M]4.���{.6����4׶����5}�U��� ytd���My4���j{ ��'o��֘q����T
�`��H���%I��9�;��7���q-W0��;~|G^�s9�s���sv�����؇��r��­�̄�t��޴۳!��[�U��b�y�"+&����k8y9�L7��r9�B�Vk����6����iC�m(�����7�^GQn��@�+kF(3!��J�����XV�����Տ#>�x�\�*������y�?�.�D��r�@�@0�"J#����*Ս8.�b�ig%`��L+�py����ϋ7���Z��c���<�yV1 �����8�8E�oX����@bRe�F���-m�}��GF�S��ʉ(��-�b�#����P_3@��9j���>�j?3T	@|�Q6I�@�K�gF"��}4+�d���qᢋ�\o��|{&G���@�(q� c��D��%j ������9)w7D��ŒD7�فut�}�f{���I��'��m�T�A�FF$
�(�J�O���)a�J���;��Ǧ�z��Ǖ��=��Y���u��n�ΆFΆzZ`|D�[*__��in��-��L��L��3�����'�M�K�q���j��b����ņdA���w4��߾ǲ�ո�� G�	����f��,�W�bߓd��('�G�t@\^G��В��&�f�r�Q���uۊ�X�����9���-��%�h6#�tI��a��2�	���v�
�I��(�9L��|]���>	�cM�z��?%�پ�����d�;c����?rn�ڨ�{zL�F���;(��o�$��̑oq��9N�4���s���9$%qש�Y�B��b���{?��<�7��*���ļU����}�	�G�2�#k��{���k�ǧ��Ѫ̈́/	�X�V�t����x̌��-����%4�(���*�`~j��Ɗ-�z�*�֤��%����V֑�l��p�7z9��7ÿU������{~��h�U��^�~L������b�\l�����C��B�yB=5�E�����K���z���k&���8@�R�G����{&�u�,3�b�n7���e�kI7���	+3	�X/���j0�Uw�j^��ƠH���<���42�\*3� q���]���l/�!�p6Ņ+�[�a&Gm���qӆ��ǲU���ܫ�A������X)���ݙ��	�Ց��z�;�1-��e�K\
����o�p�4 xވ�L!����ܝ�=1�(�B�'#_�!�f�(2YZ��o�_��e�~/u"koŸ��z0��*{<�A�1э��u�|�{Eă�	G,m�H,��=]ȍ����}{�F�@z�{f���y�V� ���^B��v�޶^��(�a6�DC-�/+��_��|Y��8���\ty�yy�á����z��Ax�L ���oE�k�����+_��I�'�56t���ldc�9 J�	���~C���� rPq�F�[��V�����D����� �l�i��߳�����?ˋ��¿��e�oL�b�r�Ո�	�ӄ��0_M���O�o�hͧ9�$Q�=��<Q���i����s����p��Ƕ�0�
\'�oЦ�Z���+�Y=�,oƚ$�魡�;t@VP�-�/+�KA���g)Yb�.�QHg�����c����
g�Km���:Y��9�.�.��53P9x�Zϟ�kr����h��fk4S���R>���a��n���v�w#���vޖJx>_�B�0�=�j8�O(���v(�k	�y�oko2��!��|�b�zz�ɲl=��ߏ~6ե3�����y��[z_%!ü5(����L��9��J�����S�j(srw>���V$�e����������SK�ρ�Y���}#��6�&���ėo�eF��R�����?9��·U����知���7j�ng7�z��7�|)�=>��3a~:�T��K�C$�jB�yo��,~)0��
i���/���&�.�����k`.��w�RG���r5 ���)J�/�]-7D��s��(�l�k����@��J�!"�m�b�JVj\k���N܈J/��M�o#*�OF��7/o�/k�p�1Y��DP}2 �4�j�hw!@Q1�y'aղ}5�&�ؕ��i�z��+���/�kaljG�'Ejbs��Cc����a]��]�I.O��|!����L��q�2�P��|3�C�Ҧ�Ȥ��e�M������h f����X8;�X8۽h9ۍn9��Z��'e��?px��}��h(�wR��@���O�&���M ��Ii�VR�'F*�*ZJW#�N��Z]ue�2$�	��B	F1|�/Я��}3j�ѩ4j^o��M�8[����8�H���̖��E�T�|��w�W<�Ϥ�對7���l�l^�	E*��2�ô��A}V>��ѝ�b��^�B9Ό���[���i�i|���μS��������h%��{p"F�9+�D�X��Z��~T��7!��8Kk[�P���)|�V]����h?��z����ʯ��^�AD
�E�R[,fv�O�p 7^.� �)�pكM�|�{��S�� ַ�}}����w;J���=��-���l�>��x�o�"�iH���+���	����P��g��Цv��
���8��ۇ9�Y�=�Z7��{������<�d��Sz��������Zp�FÑS�x-f�a���Hif��[�:��L)��0�sP	9p?l��X���M�s�L��|�6N���Yb��I&e�L9��P�l���o՞��$<w��>ߔݮ�m��m�"��GD{�2U`B�R
З7 Ɔ� ��C�\���~��"h�d��&A���t��O����@��� :�`Gftg��-���(�?>5�\��UP6x�ce�uG�t{�(лEK[#_�ʩ�z�%�C[A ��F�퓻@7ejAz9�:�`���@��r�&Pca���Cb`dN��Z�d6���o��Kmޣ$��P8�opZ�'����X����tg�<֬���-�邋�J}�J�����]/�d��7`��y���������d��̙�Z#��Gύw�̞�O���Y|�_+����ճs��%.�AW>�x������G1�>o�(���y�5X����٦�nqZz��������`��#0�ݖ� �7(Hrz�,�������~U�� ���#�G�IskI�Q���t�!���[�H�Tg�-�0U1=�$�#J�r�)�}��yY�	$Xg,C dG�$�O4�j�v���k'r���_�f#��#͹�r3����⦐�(���o��k�G&^����ҥ9�B��"�ƛ�\D^t�Vtj%�*)K��F6E���{:/����\I��(w=��;_��Z���[�j7�?')����t���bO|�5�Qٞ �7��[�����DKa��"埙S�����ӔG�2�X�M���i�ߒ$~�R��/��-����,#A4�,(Yt��7'�ek����&2$g����K-iG�#�~�l�R	(6���U����Y+�a��/[�,c��:1#��EОoA��.G�jH�@��#���)����2���	g=���OpJv�G����-!B{Z���h�U4"��!+Ϛ'0Aǡ�f�?x$	�vL��6E�?���Mw
�!�s��w����i6�yz$�Ut�E�J�<���^B!�'��ad,��('����%�!���Hs�Ui�n6r��r)w����e��N��~�~z.�;��g��Ū�d�7'k��O�綡��K�9�Lj,��>	�>
%�:яc�f0�����
U�x�?�4�P���c0=e�l��`�(�x�b�XL��4���9�3���N��l.�c�V�Cp5�=pkl3��Z���y���[��X
WZ�����i��E�@���$��%�^T6���G���C������^�X
n�E�e����,3/�\�?��.̖���f7�è)_.�X?������Z���!���F�zU��oP��^'�UHf��ňi��L���Gև���&��+Jb{���F�}�}�D"��r�q�#��F@У&uc3��2�d�tؿ�4�8� �L�������x9I?��q�t���Zo6D#�섒��p��cQ`�V���a�6m�oBG���!�f@�G�S������IJ�|,��|�����,�V�9����k����V�M�ٴ�Z3✆�7��S?Ƨ�r*��2�n�x�l`����>I3�-	�`d^����@(2���F�9�%L0e��#��YI,��&�z�lL����&B2�0�0EʉlCkX1n�5�N�H[ڐ�/d�K!�Մ_�D��*rX�V�*�:4�B�3�,�x����߉0�n���2A3�l�>d=�����%p�E[��
q��5�u���n!��l�TٝA�Ϟ�34n��������C�j�X�����>~Ѩh��?Ǵ`K���O�G�W�� ��(�~팿�DX������Jwza����I�ⵉN".I(wݙxU�������6Eܗ��ב�s�qw��$@ٸC�&\64.��
�Z��]v�a�i��S!_�n=��E"�e@*a��Sa`��*�=��m{}5�J�%�$�������d���E�q���rC8p�D��V�
-��.�\��[�{ҋ1>�k`~�	H|�}�Ӄ����-��n�"WuB1�EdF���:%׭��B���I6���n��] �I��8���%�I�����t��q��m|6q�i�I����#9%�Lۼ�ٞ~Ĭ��"�S��4��	"&ptbE�ߌ<~cH}����\�Q���#�[�h���A��b��tD�Cn>�G��U'j��������"Wn{'��9��՞��|T�Ò!SN#uڳ���m���+�Z��S7Y_b<�y���#x�$�-DA�UI�1�*��G�g��LH��� ����׭����:����[pN
��ի��֛�FW��4�wr<$�]��f�aB�f�ס/M�Z�T)��������N~�u|UK�P8x�3��
�����K�	u�=���Ss�9�ƲSPH��U"��*��"qu�ÛD��.��P>���tD�7��&��v9���A²PV
�tz�7��9~�����d��cL��@>#+?%D�� U��'�h|�C���(W$N��؏G[�2��+l�vtA��$��(�U�=��v���qr]'���E}FpZ�,�>�HW�/q'-n�WSy�O�u���+��ͮ;�&-n{�Z�Y��@NuadE�K�&MK>��	,3sj^ a����t����T���TPl,P��6睲06�Mw�4Q�N�E�+��S$������,h���I���1����4vƍ1�I�k��&S��gi���:��b����p
[�O�aWR'���GE���u�|1'���D�����-��>X=hz
z76���u�2�!JV-�ҟy6�\�k�{��>U�P9��������w�lf\���(��@� 	�.gh��l�;�hԦu��zǝj�O��b������V7�r�k"iN�ױ
�\z���O}���0/��:���^�pt9/;n#��
��Z�B�Z��2;�|]�-X��l�j/WY&ʂ�����_��Z����c4��Me!�sƸ7��[U��|�v�4�],�G��fK�K�Z��DPyaD���C{8!���)���XI�f�]��*w��Y�J��A��2���n�_�	9 �֯�I�G�!�Alr���
�D���m�H?�`��VOzB0��Q�/���=\���h���	�����5�r��i��1�dX�	��X4�hR[P�X���K���1<����Z�M�o����k6�i�3��:RV|C����hkX ��E��">EN[8f40P�IڅR��� m��N�t�I�ַݱZ� 1im��,?~Q��i6W�'ʟ���UGT����5W����?jXAC����z�e�#?�t�$��Tu
3L��]�ӳØ�đ�����*�&��>t;�w���E�V�B��OV\���pm= ()�D���aha�?~�O��5�j��h�;"m|%��V=�d�a&~S-�t��np�;�6�啸���M0�5
}CU8��-V�dO�jԂw�i68��h�� `}���%Q�V�7�W#,m���-Nx9����7��_{�!��r��b]Dx��^�m���Q�N�7m�64�%% �`L\��^����6�O��|�|�`��~�Fڰ�]9��#���pez������s<Wc9�5�j{����b�I��q�ᖙM`:a&1�y7W��M�V
�#W�5�+E<(I֏P-��s���������	���Ӓ ���or57�4�X��[$��4�3����-���ؙ�9x�nҼ�?�2Jly�۠��U�H`퐡�/�i(Z�D�C^�#G��VGD�
~R�`(��h>H��Gފ�K�7g&��}�f�&Ĵ�K�@�s��ܟ�su��=���@<ƪF5J��\�l�@�y���_/}w�����l����	8B�Y���A<��c9�+�>6L�.��l'��w����������?�[{n�8��.���Ɍ����t	���+�P��6��Ԁ��U��6�--��wQ�Ź�¥�h��	[]�Q��!��݂��:a��:��Fİ6�^��U�� n��փ��@������'Z�x��p��0�j܆�N]̟����m6��7b���"�2�TG�o7�ԲH=���6>
>h̜,~��h�q������0[I!�}F��a{��=�M1��oI@��j@���7sVA���M�&_�&y��̀̍�+������30�~b�e;͞���͠.E݄�s���-�画�(�Yc}��⻜L^���N��Uxp���K%�,��=�EUPj(|'��|� W�L7/oLZY	�U����W� ��!���@`3�f�����t��\9&�zy����W��}	ṕ{�:�tO��x�|ٺ�ZS;,]��w��激W��9����)�� ��%��<� ίsR1C�C�0�o�l���@㨭��[uk�ͻ(m#y���5#R`wV	�5��Gs�=ɕ�-�#��ɝN���ފL�#�����pL"�v��'����`zwJu�j(���8��.QҒ��Ԩi�ҍ8j@�.���Plr�Y<����a�������W�]�~��æc���0����;[턉��^�Iq#Hϱ&T��˞���O���$/!���p�)���c�cl�9�қF�j�|�<$e(J{�`o 1/*�ۭ@�M�& ��e�	HBE�"$Qt��H���F ����i�W��"�7�=3G��S��:�NE���nz�~w��@���t׃�E�f	vt\H'Q�1 ~�j�`#�Oׇ�C,����l&?����I���w�����7���GkV\�����C���S]A�0�Z�ô�H.���i��I1���	���<{�ƕG�Tn0b�1?����YI���\#�;áH�9�{D3"ZX���uS��-.X{W&��C2�ч�����v�Y�տ����j	C�4��l�xq�՗	�M�诓_��Bt�4)D��Sl�cI�$̤卌�мGPđ�"�c��3�ȶB%�7cMւ?����9c0n�0�������XB ���2b{$vڟ��d����}E��a�F1 �R�ą6;�e�x�^�&��UX�	5�_��K�k� ���<��� Az����)k��!��a�K]��f��h���|�&D]N��^�9<�T���{w�+��R���R������/G�}LD�V��"T��a�<�M���륹�-����^{~`j���P;������8�i���������, X�B�1c|���%C�Ó�57���Æ���PX�F��E��F�]]|����4��:O��Ĕ)���d�n��S(��װ�,��o-	��n���O06{L/V����}� ���#��=�1)3��m�o3�ۜ����z]MkP�y���m�m4v�j��{*�	��:r�o���s�U��B�x��y�l��rs���r��iı�G)d%����5ԅ��ޏ�Z��K��:�JN�UN��O��)M�#�j�)K�9�1�n�T��v�L�VC���޴��'�'�6�����K����J����Y&-S��Z����(~w��}�1K���|D���h�l�'1���BH�����\x�qd��A͇�.�)�!�p<����1uqŢ�V�\^u�̊��ȜF�Q��S��ӈ)X�Q�@f��tN�=A��[��Sc/���o5��6�7���f���;4����.�:Fq&,FH횧>�ƾD
�����$iب�������ʝ��B�B&C&�)����-`�?�Ex��4�<�MI�_�,fk���L���aEQ ��.���u���^�=�bO	҇Kca����y�9Q^긄Y�qS�B�5�
����%`Ru��P�A���ӽ��0ܓ	ϡa
��ʐ��D�������HV�?�_�B-(��;�]$!�B>!��Η������6�����Jx7�Wǘ�y;�"���²�� >���3i����۷
+f�L�zdC��;�w=ipw��-|�zM����+��7!���N,�-�� �_޲�����D^���,��A䜘y��B %�a��v�	#f.@�	^VJ!=�.Z�j��d�Go8r�&�'��y�9�a�2��zȊ�g/]���;K"�Wų5�D���ȫBb�
nӥ�jg�����m�֮qr^��Pù���}|51�߱cPIji�F*�Y%�  �Ae��]�vI��S�
���u���>�B�
����8kA2��C�����{����yBN�WT��T�.E���!�.��mE��[�C�I��K��M�ƪә6H�Ч���*h\(�İ�<�����}B���}��ʮ+�IԘ �a��匞�{8>�[rN�����v��Tj��Uu��J���A��{:y�,�l`K��|j]_!�_��]\�{����|������{��9q/I��+��(7�v>�Yb�}ɬpUj�{~;�"L�8��bd|%�r��|�S�:/���o���.#���|±��[yG^��ѣ ������ *���%hߛxL��O~����
j�>���VW��acA	RC z�����>4�~v-"U.�jt����E���	��I_�� �Y���~�$�:JY��U����l�~${�\�7�I�߼�1�ߥ����gx,r�3���A@@�J֚�M�P�s7$�T*4�V�lL�anD��	�:=�w���?%�)�*���NT��T�gPr���>�C~���_g�/����V#'���i	B��ޖ�oI���k��ѱ�lM�`��*�q��+�K܋�>a�%,����+�%+_`LT1��  �����ݪ�yE��
�V�,t�e��kV�L(�
�n�]�����"��;����s�gT���\bc��5�K�c�Z"�v���0G3 {��~��R�"�r���IG��aٿSձT��ƨ��!������IG?�N�~{������%�f�K4�Ba��s�S�i�ҭ��1�޲q��3BCV��"a�7��*��^P�G����3��'2ka���cעIy�?"q0V"q �K21�_���e��˙�x*l�b)-TK��U�����;AN�-؜�����4�{�R�Z1K�L] �A+FdL���݊+�����B�);A��؜K��X�A�T��!��f�$oe�D��6O'Z��q:�֝�� �v��=r��N6d���(m�������h^�3^d^E�>����ُ����a:\t�lx6ɞ4�#�����2X��0�Ib�}Y�&|����e^M'��6�|�K.���C������&k��cG ���ʠ@6���0�~E���9��ɭlﹶ�Q��z���{�v휜�[h��H��=Ð."�G�G���qlX��w����+`�����u6�I�\��	6�*�ͪl{�mT���Ĉ,�n_�!��R-���=zS �E��B)�w�QȽf��d�QQ�^IH�ڣi����Ѥ�1u�1�_�P1���5�O�~̹ �f�i?6dx���F��e���R������\���X���������w�1�� 4��h��Q�ݧN��c\)���naa�9�Q���wY^¤ȟzǛ���Ib{�����MK����)AT]�b-�F���byn��R�j����b��sq�vA���psiL��R���#��/w���p(mZ��|G��@b�Ѥܔ������	�>MV�ϵ�_=B�wA0��^�.A���s�ՄI��_Q��C��lI�79�X	Jo���o��bMJ��b?8c�a�s�QC����ޓ�B���v5�)�Vf��^-Đds[TE�=�_o�>��кl֧u�V�+�\چ�����5$�W���Sݝuئ��#7H��U���o�O/����D��c-�����]����cy������~Z��bry�z����H���͘E�
k/�-~��'����5�)�f�R�$�0~Y5c�ƿl���".��o�bg��e@9��.�-�%
��b�q�171Q�/Z[%?잪�(��a��˿^�"�O>��Hf5�M֡�XW�/�!N��Ŵ�*����^p5y47�r)�7�����^�<%�3'���P���<�"����3?�`ʸyT��� �1}ܬ<	�P5��f&��R���(X�a23"�Fgc3����Jx�j�I���$kG�s)Z<��v�R�P����
� ��P^�T7����r�~�|ʑ}�FkZko�%��v�:r*;�j��
	oR���˶���� ��G�����:^���6���;��Ǎ���{Վ��"�5�ޓM��_3e��B+����W��:�:gVXY�n��H�q�ͤ�7�J����֛����e����w_.7Og��gɆ6����(/75��t9uSﾔ��,�&�sD)���+��7��8N8+Rп��*)0j#���'<��'\�W
��L����䲸����>�M�TY�1N� :��#/e)P�d����ē�$'1������K�vj?aS�¶8T�����3x�d����Of���R7��y�z|s����!rb>�L }f9����D��q�m�����p YU�
+�1�&$�s��ye�R�FFo��f0.ПN/�r~�II9�+C�Ѝf&V�ޝ�[�Gw��d��+[#G�B�����m{���[@V��&t��p�i�����M����9��>�_&4�<�i7���w^�QM����{[�u��l7�1��C/~ĉ���P����{�e�����k;Q�	� V��U<��V�U�K���1>yn&��ǢI������j=������T��z��r��[�T�������7��h�C��$LI$bMz���Oi�E?NBa�Z`�1�.j����k����,oir69�a�J4ÉZ�;^�FJ������$,}�A ِ���I��=���=�+7����t{��Jp�A�L�ԛ)-R.���f�<�g�*�<�>�k��	�Cھ�i�L��g�KZ�ć4k��%�C�kRʐYpA坓8�Xx4��X�ؕ���'Eq�<�2ei��6* �CI_�&
�;������j��mȑi�W۱���F	.� ���%^��us�~�P��?Q��������"��'0�S��1ȖMY��P[��)�z�F$NT�	����¿}׻��ɺѽџ�0�G������t���w]�Jk�~+n��6��y}'�X5���x;���"��ݐY:+�Nc�֨RK��V���gˏ�i����[H/�@!�"�k,�f��.�i+���3��TsF����!V%ͷ������8����֑��$2����b2�����qE_8 6t�X���F���P���R֔5����)aǢb�#�'�i��q���ȣ������%:!��[���-����ۙ-�� �V�,Nv��)V�ޗAsJl��ah7� ��*�� E<\�S���j�#���|��?�b�"�� $%�L���qz���B�I���� Ӌ���9�Q�b�Ud8I2~)`�����A���F���PX������DUa�`�\�"]���:d�~5�J�����Y?�'��vAp6L{��#r�����Z����y(7�/�_H�n^R����B��ս�G��4���h����7�v�`-m���ʓ#����>�n�>�K���T!�٦=T*\}4�K�{��5�ϼeu�pᄥ��g.�@��Қ|���n�m��;��ۿ(���3�=�8�8`���H=f���$D�a�,!z>���9�0f���'Ո���ʩ2<�N:/[���ܙ�����L�X\Sxt�svb�}+o�A9��{��!̾X5��!2�AI��u4y�i�A���f^��-��˺}�;4x;���L�sPN��*R�!�Y�N��H���"�r��bR~����ŏ��e[�&��\�/�|�x�4nͺx=t�o�~#�+4��ՠ�f�����|�5�&n�E7}0a0/��~c��� *�%-2�/��1�JX\.���N��*-؈w� ��a�Rf�����O�b�����zgV����e�]�F����'?�ܓU�b��t�=���H�;l���-0j�-�%�s��#l`vLg�@V�5�_'�9�DH��"�~�k�����F^�O��!����N�F�T�B��a ��Y�]_�DI�]	��˜f��R2]�[�By�����m?�^�p��
����['-.���3*�P��S� 	���R�K��KE��vʚD#ԞV|�P�L�[e��b����Q�W��#R����c����5Jy`����D���>xCL,��D횿�,5V�,�u����W$s,��LM�<���i�ڵ�E�s-��W6ԛ�}I[Q���$��[��r���I� '{�O;��@vt�%<֍7�~�=��y&�,ޯ=y�8i�c��|�*��v���xh�i��tj��ϱ`�1,8j!R����=+�	 r�r?0�t�T���9ͩ�h��)!?�|���N�+��
áz<���9\ڋ5b�*�"㖈�n���i�F�lrUU�Ú�m
N�xW����(�L�A���'���G���Z��^ �c�r�Fđ��a�qo%�(M�29� ��@`�kǑ㿨�-��سȬ�ٻ�ة�Zn6kB���]�Dh�}
�b�A2ڨl�_�E!f�}dp����p��:�8-��k�7�ӓ(��&$@'��� ��f��@/]wO�b��9/_��7����褲��+ݏ�m�jFl��(nƺoŞQ���iܳ�0��F'ֹ�d�k�Qz��d���Y��rܓ�2yF�r�/����.Y���-��s��b����lQ������I�B���VY)yܺ�2�z;�l���A1��b�����y[9q�]Iɖ:�r��p�V�!��{�m� ��ʍ`��o�Z2��=ɚF��"��P�	�����ѠG�zc���4�0z6b�H��S��'0u��˷"��"�Wexw���^c�qv���Ub��r$���+�Z�c�L�	��4Jj�z�^�	�C��&�e���f�ʘk���Ѧ`".	����l����R6&t��fC~0f��o�D7:x����~|���BO:�F^o0�<�_���Y[��3ie<�c�U��7+Ҡ3f��1������5g�{2��i;��"�;��g��oT��I���~y�W�i4����e�FM�L�.T{�
�/R��Yߤ�u���l��_��'��bq}��NQ`�E�"����n�O	��������,<?���@�l���[Ec�?�0�+_r�۞�3��'���~�n�NQs�(�~�=�ݰ���]���l�� ����+����z#-iJ��2�lq�\���z
]�?�5�?�5�"?OА��^q�_ݯ�Ԭ���/6������'c����:'o��y_O�X�<o���p^�~
��`g�Ý/���P�/��"#_U��+i��B���0q+�-ȩѾ5�"���Uw+���ĬO�5�R%�Ms/|z�<y����:lp]U
]�02/y��Of]G ����_�\����on
�C��βCs|OphX�o��3sI�}>�D�i6�T��#V��}�e��[Xxqʎ�cB���ƮN��ʹ���#��pv���^`c,��t1g��Fw����B�}���7��X! b�w1����З��"���K�.���ѳٓz��ꩇO?���W�97|wL�������L3�9�df@�KIi;�T��DbhՈ����It/9\/�i5��{?�a'��3�}���x�g����ySBw<ƺh�6�e2��lu������B�r����z
���o�,�\�jI#,>k��{��Z��^�?�^��� ���YOj>��@�o/슡�Q��[�d�����q���k�F៻���
�~}ŧ.��X,Z	\l�;�gÌ9g�w� �К:��p�Շc�D�ɈNQ��/2zt�<���\����g%��.'P��&�Z(���e��B�.��P��J��z^�#9�ٗ�X�F��nr��_���ȝ�#d������g��}�`�~&u�,��LU� �������<e�,�cnA'�����֓����E���V
K�E��*g3�+���
��ƒ��3��sfS�\�#��b�bך�b�]�:�ɶ�<�3�l����1�o��ԝ+��z3��B-��;���r-�T[S鍓�&VL0D�n~��C��WG���6�R�k+!�]����%Q���AicK�R���zc=aNGf5���Ga?���YgȐOά�cH����0)c�;�}.;������(r��$�����H�TOK���HͭH�����B��P����"���@�D �R7A��6�fk-��<�kԈNx�W%��+��8]�-��r��2W�11�UW��]�&��D�}!�W�P�0��z]r�"S���w}C�xT%
�x�̷�`l����r�Uq�Jm �N�e����>�z��o���e~�@�Y_�}�$�a����E->�۽@+��t�O�Z�C�E�&�}F'y[���*� ?�E���(��
^R�X#����6WK�_� �Q�a
6�!
��Q���������}�����f�'���N�ȇ3�j+٨�g�S�"����
�["a�ﱼ!:~�6�>�e��e����H���3R��Je|<r�f�\��򯽏X��1��f�b¸دyI��"Kp5�)4أ#��
~x-;������FY�>�Q�N��b~1 �Օ���{,�r��\`�|�|�K*#$NA����b��=�Du~�O�6;��� �� 0��w݌��u�����a5@�z���
3[�w R��wS��7��+⩘����=����߾n�0���$M0w����UD�=�]�Kv)��n�.�rA��.����;������;_v?���9��;�̨/S��2a��N;��z..���C�_!����ǧ�����$�*��qjg� #�t��f�M���1�͞S�%Rl,2C�7&��T�8JU������kt��i�� �$ U�0��s�L+���p�_o�&�
�U��Y� �	jRf�m�Lu�w6̴C����ӱ�_8cM�8c�X�ZT��U�췇hd���6S}���~Ȝ(�}.���':#�,|(3
����h���k�vyDu��c���ݙ˓OC�-���O-Dd�5 �
ss�hvt5�����iV�$T+����|���B�}����R� h�hi�t��l�y�KvM����Bf��G� ֎S��o|���r� ��m����u\�]%�M�GZ�~%��}�af��\��1Հ>D#��WR>����9�'�'��e'	')�Z�.`/;Rat��)�Q�iE���KS�)_3`�dv������ �i�F�w&�G%{�?���K��Y�%��g.>�t�����G��u�h��&LCng�oo?�k�~ٌ��8����m��p��_<f���U_��vd�}�HOq���z���B���;�T�,��3�x\f�o�
~�W�pd�JI�V��ԞisT�媨���L���t�ͺ�@7<�&M�Q�6�
+�?���w	㝄-
���n`��Rb��[����]�v-��X�XXF����9Y f��x,�7Waʱ����Ae/h��P>;��8����C�%@U]���T���/���2*��1+#��A��zfp�1����(��= ��Av�:MKz�/x��F|��B�:ɲ:9<9�s�AX����B�z<�s#�sHb �`����Es�p!�+�[M��&���3�No� X�/��N��j9�V��Y��+aA�ġն���ϛ��{�M�^c1���_��M���)wLU�6ì�u�$:�w���y��"��1&�\	܋r�w���e̱���a�2�TŢ��r���Z��z�lZ6����I���2��"�������i��}W?����S}���I�iq��>�`�z}�����L��)�U;���4�Ҁ;�����������J�`]*����!�bk�T�>|�����/�PIw�Z'	}�#����C�HMރ01����blʃ����R�����&"���,�gU���%��c/\�J��11^jL���BW�Z�� <�޼�PO^+���+1�����@C�{��=�� a�d��
���jm�'����U޿{�&H0�G��J@��m���T�m�+���Պ���u�t���"۶���J2$��r�K�N���d�,������P0��kǚ�0֕FO̩|%��U�+/�WzoA�4l��UL��5)	�Mn*�LH���ʾ�C9� /�JK$���g ,w�K���v}�>T���+��yQ�	O��\��b�A 0��l�J׈G�����,)���A`5�F���F��$��]���ۢ�LE�E8�E[ˇ�����������ӸpF1�D��ݙ�G�b��JG�oa S����}�O
}d�(�>�h�WG��OT�Xi-_���pg���ϔn�ۮN�7ߤ
�bk���JH$������nz�B��{��C;t�y��{���8|�Ghrt:�3�3g�(ӕxM�T�>���vYwG��N��������4ї�xG�P��N�4C�c��)e[Z2s�R�T����zY�7���e�������[P����G�rɵt���-A`:�v�RC,Ep�-vj����P���k410r5�bq�P�ܽq�7iJ�q���,�H�m�[������e�o�:�_�"LMPAa"�����Ù��;�'� ���;�Kb���㳭���L��V�_�7�*��p�53<	G5�e�w]��& �@��������u���
����z3Yp�$�-����L��]�cHd/T۲����㐤�2�S
����+<�E*@C�N�⣓��
9��6;0��MRΗ^��lx����˝M�t������~]�`�S]��\ьC���I �� y��c��j�ꀙ:�@D�O�fN�|�s$���8�a��T�e5�*K�g���P��E)]�ċ{t�&W�<�d�o{Y��A�
�������v���RD��&�X�I��;�p��[�O�����Kj{6�����q���2=����A��c�� jB���Y�dfk��z�WO�XEAf~��^t�9���jY�1��v7�)�hOrl�U6�T�����O@�w౾�pm�c����wU���Amv�`h7��:v�^|�r�|%3��OF�/�(
N�q�}j`�EQ�I��������!4 c��;�SfviG7�NVϱPf&+q���L���}�Ꭓ���� �
�
�%>y3�.QvarE������[ܪ��W�6����Hk?�T��f������s�|�H����8}�"���°|u�V~&P��p<l��>��(:J��&�؁H;>�y÷?@���3����J[�!ω1�e"\���72s�MW�[,��QsK&�k���QV���<�&��1ہ�Q��Zr	��|�x�����t\7A�F0�+jbI9���5�|����P��03���ќO�?��P��~9i:l;�+���m�WbfYxJ���������R ��� ���܆r�܍5>Q��csAG����-�H15�˥*��x;E�2Q	q}�)2Y����ݰo�j�p8��ڊ���G�Z����k>WW��M��4DᦉR/�OP�g��<�k��L�'Cߏ�����7������Í�`����lP�����mR��O2��Z�ю:�'�%�/�J�~g���z�7�z�G&9_�M��<�iH����.()U� �R].�RY�v��4�<�ys�囊�S,p\�}�\�� ��-�O�����Hڊ~�zr���y��xc�������Y�<�d���c/KȨŕA#����H>1t� ��)�D5�R��(����4*	�Ag9�ƦMOy(G���M�h��7��yΖ���T��'�����`����f�lw�C�_7�r���"��m�}PLaH�c�����
��uJ�,�Sh�J�Z~ZM�r�G!�۟�{H�����Ɠ��L�ʵ`ar㆞�	ÄȤ�I�p�L`�`*��AW�N�
���R���T���8�q3#LXE?�qFΡ�{��sL����f@ȍԍ̨�{��NB��u�$4�' ���d�L �"��(C;�y@>��0 ,��/D��"c����=!1�����
}L��j�������H@���_��ᨂ�Q>�
r��7�t�X�N"dd��;�x�9��d����ţ��s�A��Pb����;�q?!���+b=|~���V��u�i�T�	V=^jI�A���E�gfIo�Aȴ�1F֮x
�;�E=�y�Xά ����1;G�8)�u2$��ҡ}�X����3����v#~C��G��^�m�\ tw �%��7�������*!2�߾>/ea�z�"?��P���]�%4ݐ��C�ç4�� ���M_���~�e ��u{B�!dnzA�����{��PY{>Vw�/��oI���?�����hFSn"u�'x/Ǉ�������	���אF��,Ǆ��o̽�a45�S��sB�����;�':���-��Ԟ�� �� �gJ���e�o��RV��dւR04rQ܄����年Y�[�Ũ$*�Z�ï�~�/�v������!������3��F�_:�_�I���Jc�X���F��&�o,��h�M��f�Dt(�_��Ԅ��T#�k�ih[hk�!z�O,�̱'3��Z��=M]��~�1�1HTZ��#�B�|���!�D��:T{�oV�v�f���W��~E .�=W���Ȫ�/��V�V���M��ܓ���[�<B���w���?�����x���C��e6P�cEa�N���]�v��j��T,����D���EӬz	���Ď�L�۫E�J=1Y|i ���7����IF��}!���f4���@��L9d����2<���Z���}�P���(j�lp�!�e�z+fStS(!`OV�}�c�q�:Ҽp����.!:|��n$C=l�|����1��ɥ��{��8g���1?���S�U���B lv�&����N5�������;H��|�`�s| ������(�B�&)�3=đd��q�)�'}�ѓZZa��(��&��S0���wn�(�ފhP��k����t1E�P��H$�5�Pi����6����.{u���7E��4r���{�P;~

�S8[	T������=����{�j�/t]���'��mB�h�Y&;�L���u������4o7D�s35I��_�- <���씥���� ��S1z�hT�[ڀ�AW��$�c�a �s�b�bvu B�g��P,ȸ=����������ق����*���y�1E?��4~f���aJ�h��cʬ�r���VN0���>+�7�@t�>*��Ia��>);��3�[BE���k�U0������, .���>�}W4:>���TI����ތ~h�PEv�����1@�ȶ��eF�_	��7�bT;��]�O�5���O�Q���9,��um�+ �g��(*�$�~�2�l��I�b���R�eocHx(E�C|�V:\�Q5������|$���-*	d+�ͤ#�%��[����u�e�?�2��ƪ%*�Ϫ�������F4��Ŏ���-��Q_w�?��w߂���)��{"�xՁ�^�����.k%����ɪ�aB�2~��h2�t-$�� m}���n�q+:���2�|��FAo ��K�Xq�	���R���a�T*>�wX�"CY(]J�Sx��y}�	�Cf��k��X@?X%��wؔ�za��� ���] 6n��b��T�<{5�~�\W�o0��[�4u�F�����g!V��H__F�T��C����ꋦh/�v@zGJ���4����Fş��ʑ%Rp%��Aܕ��P��F�3�P����������E+2(,�jڏ@p�;�V��gB]7�>�	`BH;Z��&D5C��IQ:|�(ln���h��#**�@��J�6Wc��sאC�-��GJ2���A�"7�CҢ�������O{#�6�t�.i�2����Z�/���O�4 ���C��0`��^�]Ŏn&~���Ʈ8��³�=WS��W7�R*���;���P��nMn����?wK�c��/H���4[��u3i�ڎ���(�bb�]�]>�6�y�Q�ރa+f����A��nn�f���jG������;c�࿶֋I�H?���z�Dej0��Y�Rq�=�b�\�{����>;�%kH��J9�'
�����@�D4�o��uEw�'2��|���;?Y��נd�;J���L{?i����v��
�ސ�+��Cb��y��U��5�M�x��� O�.�x��{�:��`�\����B����m����
>��ˬ@�N;>���+o�[L6�l�y���a�d�W[�cc��b�� � Z��Lv+�v>�c��o�iр*�w���o��s8�%�u��2jN �e:o|��F#�[�M��38�x��?��B��sS$�(���+��j_n7�5��#�Ør�����@6�"$(%�qU^Q��R���/����w�`��D)j6��^e5���z���� �|�t���g�|ې�䧕�Ƣ�D/�������1A�c&\�K��b��h�4���(_�i}��Ϣ�C	���ѥ# �[���Z��:�4�s7{%�1�l�ο,���Ft6���Vp�^��Ě���������0�0j��*$"��v�{� #*s��o>y���]�L�tB0x��8�F��҇���~�¨��]t��F;�;cj�&�h��jh�/"U8'�h7�����\yv������݇�=���s��0�S��R��"e�|��V��*.��'�b���T��ͤ����+i��^�BrN�Q�j4�����kc�%�F,b����#�S5x�aM�����5bF�0��`~m,�b1 o�SM�q�ii1��b6nN׍n�6��_�����Q#^������K-�k]a�9�H6:#A�5��PM)���(�%Xoy)����{����X	�f8�;\h�v:������߄[W�K�[��]����b9��@%�H�>"��}��y�)�
�*B�=G���uc�����*�J\�?g��/w�N��6�2�,��^LHV1ᎎK�C�6�(~Z�op���ȥ�n���G���yJ�nCH")�t_�1yd|n	�|�
GmP�#o��H�1|���ȝ� �wP��l7\�*We�J��L����.�z.���J�q��h��=�z�]���Z�������� f��>Lِ���V��<�������j�=��h�
7�~�W'�=���j�1;x�BqE�ϥ5�������v/�ďF��n��c����[�[ v*�5��mF]B�'s��r�������!A������ۥ��~�c��4����r��4=���ȋ�_w�u��2I���l����K(b�,e?�FuQ��\��,�3�Kh{�#��������"���g8�'�pR��U`�p�E���y��S�:�����D���/`���v������W�2��b�<�`�eW�v%��sկ���[�%Wg��_o�o���p��w�t(��6�%+,q�_��#8��K�@���}ʌ}���3���l��jr|r�ҔT<c�U�X��6'��e�<oi	��8D;
��5�J��P��'x�{�V��l���8Y�j�ݟkk�I��1ic�'�ߊ�N���Bl"�>�+�ބ+Q�~2��:!�J�\v��L0M�.$[Czs���4�v����:`�6̜�i���z�r�j�bB���3�>���ȥ8Qi$��&�|�3�r��Řk����i��G#*64FG�cXV����e*! p���J������q���%ᠪ�?�W��>L�7f�Q�3l¨�}�m����(��;��۞�[_��ϑ�u�&�)�FT�0�)4�W�a���"�)+_��|����4��
k�q��L�^�-�ޘU�Z��tm���f�]ܠ@y+r����j;��k�}�.Z��	�j[�gٱ�V����m4�X�!Y����f���a�>��D|�s��CWڮ)�X�������*{�mxH."^c*uj#>��^�ۡdM]�t�h��i2����l�$b3$$b���d�J��X-:�΢�� !o7���4���R<��*T����	Sky})�ƨ����E̬rI�=YP����ݶ!�iw�˵`�E�-�z~�#��\�4������|�����=����b��=�1����E��ues|wJ�Jm&����c��̔0��� ��	|�ľ��)B�+���h^ĩ�3S`��oF���u��t�6Wl��/������4���)��o?T�ta|3��
��[�7&��Ə�O��ȂG����],7�����O��TR�7�Tg<CL{�w�0�sk�ӏ��U~��F²5[���l-�U���^��%��;-�j�?���7ޠ��|s��ʒ;�BDA��������^/�?7Fݞb���Ų���e��L�y�:�q�|�|p�x>����1	��jo���M}��_M�-wF�Yb�I�kP��,/�!���V]��q�����#�E�����f'�y�;�.OA��6,H�=��;AGI���X�z<���W��-��=�W�""�L�i,<Nw7=ASamC�(0�Pjr҇~�����ӥw�O�	����&'7<�;0N�X����d�ȕ|�n|����2M�p��e1A��uwB�*3��OW���EswvW]��"�m�����Ģ�Wʘ��d\�lQ��k����X�B~>�y�K�P^��^�Ez�!��T��19��Cv<��(#�%Լnm��9������j���?�4JЁ���V�.��5A��uF}x{d�ӾAfJB�R�-9��>�Ä��~w�o����Nb��%�?�,��Y����<c[M���[�!�NY�a{���G�l�?j�L/�xM��d��6��[�M����_��'A�l���w���u-Ҷ[צS����м���st�e:���	䍺-5i5�F�6�쟗���]�9�u���,�����C/�,�����"��k�u�Y�"Ǎa*8�T	
�h>M�O�1f~Y��4�a���fWD�)� �2�3�XG�>f^�ۯkp���Ţa��r�N0庝�d�r��K[ɢ�y�����,i�s�M��#w�耘���J�|�pB�_���~%�/���h5�������-�O
�U�����ʳ��r�a��o�>��[��@u�n�� �X�.'�*bӼ�nlt��x�PI��Iޓ}�݃\�Z�j�7>w�M5�7I��/�ꉪ�_��R%��Ϲ=�QK�V�T�����;f�?����+�eg�Ŗƾ���|Ì��eG����]��b������J�&$��˝����֥@݇���6�?Sn^�ϖխn����^e6uz��QB�\���MJ���yϰ��r�]�۳��
��+Go/C���&q��Ǉ�҅�����<�"7��P�ϫ� �)��{L̲V$h�Hk�O޷���S��V���am�V�5�g���n�i�*�}�0&���Q��O�J#s�����)i
����\�]����ݳ&i�ӄ"P���ũw{�`X�p~�6j��`�HT��O:W�0q�}r�O��"����9���8ゼ,�_T��"}�p�
��Vl��#w���_
[,Mc��wJ�P94
� �_����)�p3�E}��t~B���9��u1�Wי�0�J̑�ZH���<��_��E�x۹�G	}��hq�h
{<c/H�͌Y]�D-vGYor��H[���mO=շ�"}�'�5��>N>b{�v��^�zMd(t�^�|=��&����:`�����	�R�.V����������;���y4�Z�q]�)c�^�:�k�^w�Y�~6l�~���~ ����I��ۂ���꓾�e�֕sPZ���Yr����v���Mx��nSCG/tN�ّ�Bm�Y���o�\Tj*
ߑ�P��|�������}>fGj��R��MMؙ��&�u8{��w'a�����_Kfb�DB�'�]��ZBto�%�j�����OƦ� U�c.[w����d��I���^D^�W�����nyy�#�*���&����+�ȏ�c*7�З+���B�f�ob��0y/�k��� �fأy�E�K��Ud~��@���"F��%-�K&��\N=24�T�P!��?ɒ��B��$]M�w�S�4�,l�� �Eq/�z��~%s{��\��-�y�-�.�{/�z�oY�c�,c7m϶�s�J��Qf�U�toa�Զ*|��� %�v$l�Y��Vހ��Pe�Z��}�1T��]�8�!<6m("��ͤٽ�}�9�i sY �Z���܍�-;4�^�?�͛��Eq6܍w�7�,U%�{&-.>y/[�oo���u��M�xYJ)M�Q[�AL@z���aI�NTR���J�D�A*��+��7޷}�&V��g��3v��cL{���cNc��5Z�vS屭������? -�(6��%�0Õ�*��`8��%bVR�u=����R�qU��~��v!� ����U�&s�9��	��}�)f�2sW�0�U43U�C�ޟ.�=0B^. <�ND��c_މEb�"a:򨯂�\&��qr��Pv�FZ�쬖,�'��/�� �3�yv�5kL2r�[��5�����k���x>�}?���r>�X�N�Lg�^�>J�X���5�";u��W������l�:d�;����<{<�^���c�s�'DA-1f���~��3��C�峍����qo���0G�C�z�'���;"������Q��n�A]���߷����ú��������	���JI�mQ]����޶�C��R�o�] �G�ʞt~�$��$���x��?NC?��@����
ǺDN��R�7E��EkǄ(C��ͩa�,�1�2��|e�u��I�����7��U�]٭>%r�/�x�djO�-�+�O�mg��x�<�*U��1�=_늦:�^
����KL��LH]�L�'l8���V�S.�(f���ge�N�A
�!�_����S=^
��*|0؎P��	���uU�Ƈ�锉+H=(,�0����A�şԟ�۟S=N2?�{͞�\5^_�97��K\IH����2�,Hψ꧲b3�e��ݤ��<�nʛlҟ����K؎�b��*Y�3Ǭf���<<Y(�,�8<ۖ�\�-W[/�\�X��=럯��4�>?>t.� �`�4�	^�Kon�mX�]\$��Y$�?�n˩�k>��~$��~�p$��>���gWr�*u�2�6�d��,:���9�C���\B�й33��5�v~8J���}�����ؖa�>�.o�o��X��<|#M,�h�B�i�d���������%m^���ʦ/�!�A�'��dL��J�t����I�!vV����`&ܺ��)�s%�}�b>[�/��1�>d/)(��R\*�d~��?���)?un�<�-X�۷�<�(V�U�ˢ_�&z{�ʻ�W@�<��H֒��<t?�h�I�G��ar��L����A����Jd]���O���+�MQG��Ke���ZAQ�J��^�W����֏�������OM�G%��֛u��������.�S�����&
#V�W-��V�e����;���>,�Ώ�;�{�o�����Z+~dO\�J;/w�����8!�6W��.�F.��U���k[��i�`6���Y��
�ģ�>�p�^ta�^  Kr�bG�0�1]��i;|���o�����y��voTm�_���=^=�XvS��%fJ���co�C|\4�{�e��/<'8m�{���j�^i�~;�8���v�xT���k̃��3[��ǭ��Nm���w�������S\�P�x�ʾ}s^`��|^����Wن���>bd�����THz|�v�P�:�&�U�f�*��E#�a��δ��G��᝱�(��4��
���{g��M��u-����M���ֆt�}y��n[����m�$�9G"��K�ˎo[��7sɛ�:���{X-��.;�/$�l���oq�W�x���`�(���V�]O��|�ޡ��Z������~p�t��t�#}e'�\u?>���QVGQ1�|dR��yxD�px}Wwt��{����	k\�W$�N���wM.pބG��~���m�+ �מ�x�9���؍;<�6Oc*����}�
O��UfR��Q2��jR���Z��Pox�=���1�*��Y���p]�y�����/��i<��\ŗ��Wx�Z�X��pg0a%�~�5�9���T~KN�y{}���$���8|�Ik� �>�'��Ey��Y��AL��N%$�Η��Þ%�a����Hd�m2lCt�L㾪��~�I�Z�?j2��d�ݺ��1�^t�ӽ�3>�&�ڙұ!��j�b۟I���:Vx�������u;��xl ]�[�����oW�8�gԥ�w �7��L?^vg4��,O?�f��"_ٷyw�/��x�>3Kj�0�m��la��eA���a�8�E��:��ʶ��Ƚ�G��q�삥~�ӯF������A<��L!R���Go5M��g�]�)������q9Z�|C�I��E�O�G2�+��o˛�ĳqj�a�����D��m:��F��&s>@*�~Ͱָ�~Y?�<&>=ܞ�l��eɮ�O(�ٷ�P��/�d��E�O(��0�qj�-�T��޳�EQ�wִ������$z��|���c���
_{բ2�$q{=�de	�*�B3R��k.	毓�~'N��r��WvH=;�<O?_O��r�%�|��U ����5�t���E��es�^��5�C���G��L��A�ͮ����YXq;�?>hY�{�`	�!�t�47�/t����\��V����о����lD����y�!N��+|)��Sг���ls�������|��������f�{���r�n�#U�樹�)�#1O*���/Ԥ�LȭA9G�k���v�?�4�ɖ�n�#_d�ޥ7��K�<c���
�)������ngG�h7���,`���d�,��7��oeD��cE�@FU0�wVm$��5����h��о�.B{���nh��V��䇹���.������@Hj��� ���"��M�N�cELC��Y&E�A����`�Pm�.��G<�k��	Q�ͳ맅[�u�(M��<ߜ;����i���߬�n����2�#x.����ɝ{������#�=�jV�u�,�.M/�<ȝ2�����]�;Jy����{�ط�:2]�Y�{�b�����ݧ5����.�n�~Z�|�/]��!}��U{��k����e;��S�#��J:H��L>C=�/[� ��7
/E�s�V! =^jY썡^,Ѭ^H�sXHf7X@g�݂r���������
5�V4Oa�F8����u��ډ��=`c��U�T�,_�A���^��D~�I����އQ%w�|ӷ�J�Yq�+{�d�U���mX˻�4��,r�4\ ������8}�+�)��6�C\�^�e��w	-k�g�����/4���*��|*������^X�B{��>i��p�a<h�ꡰ?�;������1��yٻ7�����vۦ�rJ�>�m�([�fō/!G�>_4����x<c���6,�n�v��HZˋ�����{����qS���C������ȡ������ �շ������Eo����Y��?Bֲ�j}�dmT~&��������r�P0|�ګx�0"xN"���6q^�p��s4gQ>����a�Snz�1�+]�N�'B�,81�LA�ai���c��_����kOL���f��!�b]�U�y��˚S�g<dtu�
�ŵ�11�D�-�6����	8���U�J��c��ί��JH��>$�@�S_Q\;k8��Vp�ni���h,�+Ğ���WF�q��0WEVV��Fg�3�͢ÈP���W;"s�K�޷]�Y�Ds�f��=߬GexqM���(U"5�~���梗�/�ƶ�h���!�˸��Y xގ�/�趺*i��x;�ײګ�yb:B�ު�|��7���W�{�V\��>A�N�n�HPjy�_(9���{��n>�~�����赲W���eo�eyh-�O{�n���(�g��J�(��w��VGg~��7&q���0�X_�ҮP����v��E~�`Xq�_�U��Ҭd:h�O_�)H���]
\��Z��S�ґ�Ud=����V"}���K�T�s� 0�W�yU]X�'X9��Mg"ҙG�1;T6�ߦ,0������o�:�"�Ww�? ���}���`P�6��Ԅ�,���s����IQ��2I526��1.��[ӊ�y�ϫ*���e�a���>�vi65��������f�S�UebH�9Q���kq$�#D���a��s��
�9�{Up��qW�"�Hm����3�������B��y����{��`ï� ?�(P�26b�S�̟5�"�i�J&���%,p�cj����E�l�1{C��OI[�۶\8��%�9�����VeP�P��/�_Ϻ/ĺV���h4±��T+r���9a���Ԣd����a������D���za����|a	U��^�`���VLU$��|A�D�r����'2�AT��E�\��l����x�,?&r��eٳ�}-�^�봋`������~��bc�ĺa�Q��љ^iݘ�<
��W��HE�)]�k\�W��n�����U$r{����WI�l =&*5E��8zi�GH�R�e�i6����������k�2au�]t�v�!}ft�
�*"�\����j;J-b/���m�(�E^�_8�ځ��B��Ù,S��?���E���Շ�$�鯞n+���n��l7�	e{`�}�eҩ>�&�U���6D���y��qjbm��qI��+��|p��;y�-,��^$�2��Q����|�QSSο�˚�WǕD��)�ɸvE���Z�����3^+�J8�a�U���9k*ģ���"��_�΍�w-s%���kd+	�Z�rM��
9�K ���E�ǔ'��~��:z���E�R�Gr��;!u=�yZb�g�I8`u��s7fQ?7��7tR�UI'�Imt$��V�?@�5@i������?���ȏ=1n@�FS����_?�Q�W�|���Axڛ��-���C�#ܲZ+���X4�h��u��V��PH7/ƕ\�E*�g��$�z���_��O�z� �e���I8"PIڠ8^�m�f�m��qг��Gz�e������� �6��L�GO���'�)���W���
 �+��q!H����C�YE�6c��V=`��$�1c�l�(�:	��K��'0�������R��/5�l�f -�a��ᛚ.�'����%rFe�2�/����?m�E�c�`8�	�ַ�!˖mj
�� z�©o�he���7����wV/�UC���T2�M�ϭ�}�qF�.����\��ah}��+%U:�x��0��(t����y9i!�֕�DW��b�`�yު\��+��?	�� 1Q;)l<�f�'����v�"<���V�G(��ɲc�hy$Ԯ�*�I��<���h���$�T��H�*��-d{F+��q�%�0Q�� ݌�ع�`#��"v*�R�u"`�W���<�ڋ��B��<P��vϸ�f'�JD���,':p�bu�>=�����c������e,�"��Dp��F��S���\(��AYL/8��*�:K�u�_g/\�,_��@�$��m�_g�_�=����R��~��N�9���3��pZV����P�/0�׊F����F:ylQ
w~	Eum\�H����'�3qW��/���@=W���1��og1ǳ�za�UՁZ��qL)�+�d�9�ǆ�@����4?�}T� ho"Bd|��j�B��N:�n,��-�E[��7otl���;)	��uT�qOS�tp�qT��,�}���9�ְ��-�K@OU��}x���L�bki��@��sԸM6��~|��ܷ�g�+wIȞ㤰��tց%`��@]����L�u�@KJ��t��͑�pq�KB��x Q�����u MG������d�7D}��A�3�`С,�����[�	��
/C������"�R�ҭ]_��G2�/���kvj���is��9 �  &��gb� ��]X�IdC�U����t���17���[�D����;y%0��A����k���3�)]�Ō��U�u5�y�1֖�1�(����Վ �W;����ص���Ҁ��Z�i|���v�H�.���O9����Md���\��`� Q�U�
�g+��X����[L�3�b,d���W�ab������U�;�6;�_:�UQ &+�f�Ct�X��T�Sk��Yx����EV[?�J��o+v���php����L�'m�k��W�����S~�@�^QEf�b��4JTe�փz�C����y>��W���c&��Q�v���Fmxy��+~�eYj��� �>��b0G6�����#$���F��,ZH�
�"6ї�<��S��эk�LFI�C"��b�w3~���,��W�۲���ׅt�p,.4:,ޜ�W��V�����u����V*D.����HH�U�:uO�䬔w�gViL~P�1+��q��|�Z�_jF@Ly�'UV�\��������e��K�ض3���;�29%t�o��э�x���ٱ���ab�v���8=��27߱gh�_�I!.�`9K&+<���٦�Gc��O��h�kܚ�RO�Qz�A_[6o3_�y�|DĻ�H7C�s�p��r/��M�&��j��$l�T H�	��R��#s���Xm��u����#�lTI�f�����C� ��-Z�J�Uʻ�aXw��]�a�m( 3*��V��m����'`)��G��U�倸~BW�BkX[�@9��@9)
g0�ӟ�u�ǰ��W�w2�q��	&Dm���An�;x(x ��i�d�/�*�Bd�U �nt�Qڐ����U��7	�:������Ŏ$ᱞ����RJm6�i[���j�7Q�9�[s�r�Y�p�jg��l�d����?��������r-��<��9ɩm9mеUT!]Uؑ����(��٭�Y	Y6�ym�5=XK�^��xlHe�:ʇ�B6�I���#�����vD옕4��M��5�65���UZ-[���]��	�UjSU��j�ZEͶF�7��?�s��y>�>�8�9'T|��j��6*4gWi�yl��T���L�{Mx6֦��h�7�AbƓ)�	fd7��E�u��
_qS�BT�|����S�#㉺!��Oo-�)(�TCwJI��ƹپ�g��]�hv/�zޒ����h��vZ��:G����lR2@�/F/5];��?h�yۮ�\\��;��߹�ut��F-4~!���z%,(�CW��t\���A��H�|�z;K�3����Z���0��:b|�����������̱w�]���0@�J�L"��R%������2F�Q���xN��	�;�$C)>����"����tM�F>�DNcB�'�NsC�>�R�ngrf^=$[(�v��z��饍v��������7�}sm@�E��f��rN��$G�$�=���}�[MYīprlB��W�{x�Y�z_���D�����s�Gl����_�ЛJk��DՋ��D��|��`�r��y�j���{^����R�!��]�Lx�n��52C��Q%��_�Iv�мz��[3S�K����&�\1�S��(�r4�W`���9T�T�c���[}���S��^c�,�zn !jq�!���F9��Ձ�Ȫ!Z�, ��p�`����L5�2?,�e�����M> C��U�[/;3���xe"`U����E�d6ebA��^P��C޾���o/���J�Lȧw�a�@Rn�b�XVݫ�*��;T��S�м[-�Ow�UO��T��h�l5ި*��JiA8y�k�S��Y�S(��Ze�N����K�ݑ_W����.9d��2/�=-��?Y����x,����弗���Y�>bF��@��L���#�kK�$�4�Kb��+_;�A,.�苅��NrT$N=$6��vϾc���&\��j-��wO���,���L��G��ӽ��ÕrR��KH�����G6������C�|��@X�9��!q�XyQ���c��;��f�|유2OdN��gOW�WX���t��*ڢ�ı��xx�3
N�����'�p	L�w?ɓ��1j ��G�Rk��RG�νO��U���|Sg����N�Euִj%��8��_�0u�,XW[eYbT��%J��ۋ��{���D��a:]Z�����l.Y�1�%z˃�#ۚ��,���Y)�<&�G?�;2��� ��3^����H�����\�#�vsd/���x)�=k�u� ���I�=�q�#�J^.�������r�h�N��Y��K�&?��F��\,�)S�#�@^ ?����q�^~�J����l:I2��Z���T�e�˫��7�_?��<�^0����7
���N��P��4��g�7]�ǥ�֫
���];h�K�Y|�q�t�{rE����&��e��,��3����wd�O�X��Ч�e�Ip�OPbm�,r� b@18�^ᮩ��[;1��߳����v�^��A��w�(�<|�٣�e�J��O9�H(jg>~D����cuq�[���$��|�magp���'�"�<���(�p}���{\�@����1��fvB�t\o��,%e�!&��YeC�湾� ��A�p������y}�7�1���	�h��h�<w%*-SX��i�h��x���)��#jg,G�;�"��kdQ�6�h +���-U-˜+V��e�j���}ٿ*��p�n�y���%R�؅<�y� ��^��"�5���b*X_~z:���SU���?ƭ������Wil��8������I��\���5җ1��xk���{�ٗP�<`b��E_�O�ǧZ|6�&ƚv jZ�ğ;"�e�N�;�VOL�˷��?�]"Hj�h>�]V����<�i�qo&,&�}�]Q6�pU��`�@�T�\�p���b*�U�����E[�:�L�排�����[k@����|1�4xq��3���_V��2�u\�A�b�Ƃ*�Gm����5��DɇQ���G�?����*�?3����!7X�����t�������u�خ#Q��K��	u��ѣ��:СO�̋w=�Cofs`MI؄�9p?�P�ޏ��I����#���{�gJsl���'g~�����<�B*Oۄ��������OB�1z{�]8�����]T�Zo\�C	,���
�8az+)B���H�ŋ�~�ZI��)�}2=ބ.�s�~ �N�ì[�"��oUx0]4ʧ����2�2/0|�#=��J*�L��l+������e�$muV�޲�n�c22#�[���Q���j %�@M�Mt/��z��.�OAНF<�T<Ͳ���W{�2y�}$A�����<��W��m7g�G����b`n~=u�kR��8��U�g�*���Q5���[�3"B���R H����ڑ���@��H�Z{S���֧��~����9�B��czw�Ќ�ԇz��m�:I���I;����w1u�t�u��˫ƌb�jŒ����a��4��T �*P��^�#����ҥt�jL$����*B�����5-�^��xZu(�e�х�6C�����}'��:bV����K�v�)6ZV��3��|Hq#l��3\wȑ=�t"�j��л���zk���;�||Yxj.T��+��/����~>~*)?������f�
�ǟi{�G�慷�2�V�Y�<�,�34��A�)��C
Ǔ :��3�A:3+E�b�a&��*k����v����&�h$������rr�n>>I��[�7K��՝���)M����@��"J����|������6e|i��>a����Ziu��=����K��$12܀정V���V�}lW�\�0�\k�'t�I��!�X���ƶ��o�9B,7�`�� �H���rhŻ����2������gB��V#����Y�����}��i1$�ֻ���|� P0q,�z�rV�5��A&2���J�r'��֪KU��t{��H�c*��<h��`~^��go%��j(I�>��Oۉ1e"Qb-�W�^o~]lË��Ľ�7��h���!wZ>��\?�,c��X�B��uI����5`�^�i�L�ʫ�ݱ�������~T���~��.���g�$	��Sw�p��+!�B��&(A����d�F�Sᢱl.�DJ��r�M_4���Wͩ䎻Z(�̼k��'�
i��4���J+J~�1oQ��r}r9��/���t3�PV�Đ�p�nz���[�a�V���RF�'ai?Y8 a�W��RK� @g�%-6�AT��������M<�~QY����R��m���SVd~����|POX�?b�Q���R�0�MB���C��q6���/���P6����FqB�}Y;�Ⱥ|���W�p�L%����l8�ԣ�r¡6́T���6����d�~���C�Z��P��$O*n#����	��O;�H�Qf�W�=��=a݋B�=$!�Շz�]�O�SAjr&�M���'�"`��_�E�O��.$"�2٨)�}]��BQ�-�u�����ܗ�:������S?.�(ZG�G��P-�m���
h+�Η��SLN�{�	�s8G�]���pC��&��p�S����hc�d@U\8�u�Q�]��7F�'�V5�����������/Β�O���������p�b�@��`-V|���z�P�����k*�H��.�5;�jq"�7�i4�z�d��t�K��w�.��y�fz�gq�yƸ��b��=�:D@���s��n�ϐ��<���
=�\�.�줻�La�;��T�h�\	Y�`Am6J:�䗂���!M�k�$g�� D�SU@j�\��"�7S��r�r9x0�׀29R���b�h�N��%ޖ�l�O�/�%�E�'���?Dn���L�g� ����NE����c�@	QO��Q��ϒ�za_N�@aE~&z�.Dg���i&�ou�����X���D=�6�rWG1��=X��vGԩ]���A3�Z�����b:��I����L8x����9��=����.��0�����������T�,�1��za=�#�9��}nv�C�̻ܠ�ٸ���S���2�d�����Q*�B@�CSM��|��$���"z�n;��W�@a�8�z��Q����>��� �R�����cŪ���9�W���b��bC��I�wɟ_Ɂ�U>���~�}�f0S��3�����?`���G5�<�qȅ��uX|8�r�.1�P!�]��[����f/�,?#j2
��/�G\�����1LĒv�~.�)���ޤ+�<�> �d�X�I��"�]o��L�Jc㖗%]�s/;�T�y �WG�p{�,��it{�s9��P|����[���i@�Q>�B	��\&��Kb��k+��'������d.�����8��;��e�2a�h>-J(���,����'�4B��A���C��xE�Q`�h ��l�k��7Qb�Od�瞷���~���ħ>���[��>U膥rA�0��cI!سV�
I�l[Bw�^"��S3s�".�9p��n(<�3n�g9���<.��MC��}�X�j]=Bjʘ�r$ĤA��B*���m�AO��`�JV�}ˀ���gA�� ����1���l��Q�:z�{�E��4�� �INŌ��'�V{�]��4U(�2��yِ=���u�-Q:FM�3��[�ݨ1׊ܿbm�(��&:&<J�צE^�B�0g)���6��V^��@kY4��E1��d�?��o�4Z�2�}�m�Ld�z�.���Y���#�&��r�W,�׋5�ц����L%E���n�Y�}�t��VeB��|J2�R���²��m�r��|6��߄�iX��j�LS�x�eAO��1Ҿ�0�I�QtoA&<��� %"$�� 2}	��PT跥�Z.��哯S��=�t���ט�����#|��+o�@�j������Kx��+�V5/�t���^�-ar�3ʛB6�-}
��a�$IK�ې[�bY��އbQϴT(�_]+�M�&�����H�X�{ [��LΎ`������P\	_ي�J�Dd��&
��뗋�mc�Z'
�RnD����a��"~tUS"}s7��bw[R���|������'��e�*���RV�bP��p)�W6�삷1-۸�跦�h	��:���רÔ��ֱAؑа@���GtM{����]��Pm����,4�4��x���JB�a+�������:��L(�SH=��_��%���S�x^���st�O�����!��,
���aM�ϛ%�VR�^	 �`B��1�$�J�p`�H�Ϥ�_���	Q��������c��;S'� �M����q�U���K�����ﵹs����g!�-�>Ŋi��Я��B���X�MY��1RQ�oj�-s�Z2-���"���6��t�u���:=z�-4�C@�t�]�YK��0�
���fP�ē�Tv��*�����uؒ�̐Ŕ�}C{`��:T�ɵO����u3�!��Ux$��)7���9`u�VyIg�s��h�L(ܜ�ö�R0 ,���������m�ͩ��ǐ�U�	-:��[?��`��S��y�>'�|f����e�t-�&�8]slp����X�T��L��DWL)���I2���u��H}�"B_��0�Oż���0 ��jw6a��!�c%�mh�<"��>�Rp�3�C�V�4�����ǅ1&��_��섐]��U����Zo��N��Y?4�p¤�F+59�U@���7Ӥ�*
�;�""���P*�����? �z�h$�� 
�Q2$�[��o�o�%�Q��E(���QM��h���T%���K���.��;�lU�o����7M��O�À<#������:��7���w��x��T��'�Y�"szb��/7Y�T� Л�5'��|�� �i^w�r�DSL啍I�qz4�����i��CFMl)��|&�րZ�z� ���}i{��*��?:\\�����Sx�:/k���g9�t��P٢���lO=:�S�<a��9|�׽��?���''���&��:[��
;����9Yv�/ #�J�/��ɁMF̩�|0��hS2P �,�I�����#�ds5�-��RA�z�&�y�Uʕ�쫙9�%AA?ԨJ?{^:"�1���P:�BW�	V?�(/�v~#��G���"v)[{BIN�3�y�����Y�=�^/�{���^eS|mt���s�(�#�r(��O�^�Pj7�D�S0a���po��1[��\�mO����Ti�C��́��'t��UJ�(�cO|g��p�R4"�U�����HQQ�#�xv"�Vb\B�{Y3U��a�s���E
V�l���ukC�V�8]>V�}ߖ�Ƿ���x��3n��L���߀��rh��b;Ъ�O��a��cZ8��c��RQ�t�����m�W�Qצ;�B�B��_�cSN��͜
-�Ep�ީ���9X�tw;ȅ��#"������i��.��I�m ����Q���Vv����)c�osd���b�*[#BV�f�l��;{�&����]5����+O�!��~��6��6Q���|UU$ա[M��P��DɩU�P{�P����Q����C�.Z6܂��@�����m����Jsj*����q�� H�0�����의�˭t��3�-��,iX������Y����#�
Ɠ3�=��{��/L�g�г�J����״�a-��x�'mW�u^[xT�ϗ�c�c*��ZD�PXe����KW��z��{�1��Q�������hSY0OS'ਲG-&�ױsD�Ȥ���Z�3�߳���n�O�h�ag�� �=�Ce0}��+�s( OЄ�2}�|��(P��"
�-G�Zӕ���/X�-�>�p��}���dB��k�I�Im�J���m�ʈ����J����6�an�P��jg$�R����Z����3�~��"��ׅgU���Ӓ���
*l�2�*x�Q���j�������k�7B�����"1���w������K��3�����Մ8��!+|��´�0��z�i*`���rrd�́�/&�HϴF�EH7*O
�/P^�g�*��ow�v�F�,��|��i�uH4�Q0�|�Q�h���5+v����{e�E�뷼/8�T��s����STUY��C1�K.����!��r��Ch2+eRA��곏{�	�"��|,!kE]��#��ɹ���[��y3��&���}�y�j��|dj^���� ��>��o.�[,�@e��[>�_��;���⧎_�J?�:�����,$�};D��!�i���D)����p6�tq����S=���o��u�z���}���߰d��맬&��r�d�:&��1���c.勉�]Q��P����%����f��k��Ő�
�:��а���n���ķ?c�vL?��X����F�����vQr�a:w(G}@��~�Z;�
Oe�WH%H[��ٛ���,0z]����e4���z�d��="*�����v� 7ب!��Z�-+]kC��q{}.��o�#̘R��yF�`�TŰ��0^�0�t��'��/6��?W��`3����׏�0�#���Z�^$�Z�3���qG$�aqv��GprE�6j;��7״K����U�$;�.�Ym�Aiyl!�H��
�K_�nH�ú����ʿ%J+\]�&�h��@C�ű�$�JY�eY�΄�V��ܜ�vO�����c���<��q�H�:�t���6Vo����_��eW�,�!��?��D�9��Ā5jd��,����EF��w����۸H��u�s�֚���7�F��b��{�\��u�T������٫��hp��W�OKv���6��0�D�ͳ�D��&9�dq8�Q���qG�D�r@�B߈�8�i\vC�)
�0O�%�@�C�F|q�G?6�3���Eb�)�VH�/�+S_'K[F�9���J����EJ7O"�o����#t�ٴ�l��ޯ�ku��*�CH'��M�T$��V7";��e��n�^Z�g����o�f��vP����� _�����]v��ME�	Z7 ���W���ĭ,d�P��I
%р�[��~���hAO��^p�5�,�8����m�r��J����!�#I�Zr\�=���,<�*�3!(�5�n�N9*g�<w+S�n�V`8��r�빆�aўS�m�A>�h�A:��唦�#�>���2V5�VZ�]:��[��G�0�U�c�BIq#&[V����h}r�kkԎӆQ���Q,G��:	�ZE�ձw��Y���1p���4�g�N��pF���|�YhY�Y=X����Xx������!���{��C��m�8e���HTY�d�ڲ�w�����+�Ų�� # n�޷��̦yɌ�"F�cZ9M�MUq�8��x#�<}�����p�ua��z�)Z��(+��OJ���v��vie���Q3�
��������5�B�V7�N�V4&I$���4!_���o���Aŧ���9�����[N���"(R��S�f�∾�?��<��jQf`b���/!����:�֗� <��u��rTCA^�Mb�||�mת�$�S���m*�W�wNP���&�����WAV��������k#�N��@����uY��E�h���Z���{�l����ɝ��S�?f2��y�������ã��l� ��+��Xvd�_J,,�[�*xj���O��)?!�*�-Ja�G�Mu��=r��V9�L�b*%B��H���7��e8��_�d9�i���O�����&Do��|<�iq��f3f!����;MY��������	�����|Qb`�d�G_���4Ʈ��wNH1v��m���$��y��m#)W�x��]�Q�h$I�C�� ��ˊ��C�&��l�Ni�V�H5[A[�,7���<�({���K�?�f�BI{�}tv m�A0���42����f+�/�~M�,� Ic��`Qe"�GOu"�*G�	N*Rw�IP��|�2d���8 �{�%�+�I��_疢�̀v���ֱ����	�@zEŌl�]몢eE^&GX%B�Z|��l���l�"�����)a�xcC����J(k���:���v���{b$��u�wB՘�U6&u�e{�/��&�_7 i̓�cp� �.�7���9����|�X�(�`��m�t���Cl���A�߭{�F�#�:��X�y4��2�ww�n�d����)���}������1̑��^;}>}�EXT#�E�,Z�FTd[׍-����W�;@�CT�!���Ȫ�������'<a,�3�[�q�6�(d��).�q��Xջ��l��~/���e!3}�EJ<I��}@"5�&��I0-�Q��5I�+�;�N�(��{�Zy<�3�WT&;�v0��ԟ��e�p:f
g�`�U�����h���Z ]���Ki=o3p�IF}�>N0�rӠRWr�Ӑ�\*�)���܉}>�zgM�6|O����̿/rN�S�f<ץ��W��U;�ټilLǎq�v�A����\��E�X��eDr��ǅ��X�jP�$U�+t� ڝp10\ۘ��E�8��jx]v}�h�E��%�95�Ib9��_]��ilznЎP�V�(�0b�T-����=�g��z_������b�o��S��V��C-48s �����1h�N����%s`��O�᫮s��<m9X��r���j�0���� �.�Z.;O1rc�G�y��a��!7k��b�h�Y�_�+��6��pnx�Hgo�3!zWX���9b�/BP����R�-�
���M� ���mK�\�~k�W���D��k}��pr������u{u�R6�h�e���y2�J�.w�\k7*��O��O-]�NŪ��A����j'��!߁N��]��05�T���� +��_=1V������pE�|���2��_�"-�T�k�ҡCd&��	p�v�&-�??8��iHs)0�[���@��r�u�^����P���5BtHߞ�I��kGa����9�&�u���ۑ�)�}���vp�p>�!��C C@��j-�WZv愠2�-+C��Xxi]�T@�u"Jԁw-��L	�шqG��L����^��ԥT��ūn�7j�<=�ZizF���[�[.��5��j�|f!~��Je�O�ɟ�'=�1�Rs���d
��0�������SVv%%>��l��8��Rz5�?�Bb����T�#6�I�R��^�&�!pC�C�,����w(~,��L�{����g��c�������W'���Y�9I���o�!�����������gm���Ղ��O ߬��Ruj�w���;�Ӕ��L[gd�J;Q��񴢛����|>��';:���Ӆ��~!�<��>��]A+�޾�N/2�I=�Hor`�>�����/�Ŏ�2(�d"A]�F�jR��{��NE�H@d�w��B��8��m+lt��:���-$R��$�:��YI�p����5��zc͗�eÔ}F�t�_[���W��t��_Ϩƭ����{R���3Q~�=hO�_��K.�!�����v�Q��q���ɩ�e�8�j[����^�������B�?� �� .��/ڰ�a����yS��&s#ͣ[�U��fv�M�_"�<G�W&��#�Znq��˯�7C!)xD��<d�uf���Zy��R�����{f�n�}Q�s�}�@nfύ��'d՗W}��\�F*�r���C�}�TF��bEٶ���=6�{8�x5sg�.p�=�P��@����쵃���)�FC����ۇ\��u��S��[��/�{{������%y�(�B>:N�>E� �>~�i���a�&�<���۵)�n��,Si)2s2����l0��S�B���X�Ķ���Ļ0��7���|����X/*r�q����&1������,nu�<d.^�ق)���m=k�&]�lH��r�*̭a���(�i4�6~e�7mci�Ik�C�4�V����8zH$�G��O9��H�hO���3[J����^��@�X۝�Y�!� �ߡ��fƻ�>�A1`΃��L�j����%T��=˱����K���T��1s���?���s_���Z?��Z�����^��=D�s�@�$�R�co%D�������&�}�>6�N�7TfY<�Q�Y��;����9S������.iO4������e,�}�Չv�ǵS]����(�h��K:;���z�c{�I�_p'��,&��8c��C�����S����
�h9kg/I�	,ce;ؗ�vT�A��;L���r+ImK��?�"�,�1J�漞y<�q�cx/%���i���S���y����^�]�L�S��<�I�����k������к���۴��h�(K�-K#�$�+�Ǣ�^�N��L@��]녙tc�����b%�-"�Y�73�Q�X*Qg%�1��y,w�<ˁ܌���������J�rd�k��͈�[�2�5H�q|�Di?�l@�T��4u��̭�c�&{�������������M�6���7e�h伭��0f�X�ea6`�w�K�A�r��wܯ�I��?��{?+|�g�)7�yq�4�3-3�X�����N��;�S�pZ�>�;�!P�-'����4��� ʝ�����ɐ�I������~[�W}�e�{#N�,w�5
��9��؏OU�-����|�s=���ƶ�/�a���k5x�g��P��U�w��[��ixZ��|$�ڼ��Ώ�b�o_�)��U%���~�$]Ӧ�}}�QL�:���h�z@3����Uo��)v̑�{v����T��&`��J��$h��]�?0�ʋ"�53�O�q'�i���y|�Ӯ(ߔ,!B�.ճ���!L�qV�m��|��Րn���/�x����7��S�,i���Bx[��f��
7�IB����=D1!]_"�}	� ǰ�,��a�����V�)�u�1Q8�\�t�������
��;d��ț�J���$mu�	���a�?&��k�iy��F,=d������2��,D#��~��j���?[���o�vo���Z��no�����A��#����U��5���_��C����A��{�!V�������>m������FzI4��2�D���T@%0-��O�U����j��ֿGm�5a��K��ռ�y%I����"�p�-���־���=S��1I�RN]�ɻ?z���M��'��z��}��ߡ���#��-�a���"��O����v�M�ݥN!Rò0Nك��������"�ez2ck9H*(��׌V�.�����b�Zt��|\~>�[�f"�����(����lF�J�ĖC\;7\�rt�є��+�-��5�T���p >�:��ѱ��v�v(@���E�j��l!��Gp9͋Z����6B ���j��9���X�vv� ���U�݈!��Zn�����Z��)j�Ts�_B��cJ#��	���N�55͍J/�*�<�WF���^2�)s4
L�Bv=�L���{��P�D({\�ln|c�.d�{k�_����fM�%:D��ꍽ3c�6#����ƛ�Akï��Wsj
��8�}���#��A���;w��v雲r�4��"�3(�?�<3�6��-:��d�ӷ�%y��,�sՓ��_:�Y�JJ�@%�(���݌W~�~N-3Gl�W2ݫd����}6�5�����p�1��15��W��?�F
�������<Zl��wsZa���Jw���>ӵ��-����G�~��k�N	�b����p��fs�}�kv�i5�B�PѼ�ey�@��u�E�Rud$��u���o�~��:� IZ�\�0�+�/6���_!:.����GŢ�E��c߲��k�'��@�:�W����qy�z�	&k ˰��J��1d�o8���"�F���fCP_F}�p:Hv����nNk,U����ǫ{�����+J�R����>g-�}K�Ԇ�(U��B�t`_�e-���X�
��m�qS����ey��/�޽���������U�g@�BH��z�n�.:�5��&���	�L��D�fm��qc�ȼw����"�|����?�6��Fy�&r�v=�T��`e Sa(SF8�ٓ�O�OI�v9T?��I⺿����/l���E��j�oaG�R�w�����;�p޲���Z��X٨��P�D�F�h��d�> �ׂkb?�|�I�\@�����p�e��j��Zzq�	ʋ���V�����X��q�ǕP߂:�+�60�5���6�υ��߻w����(����R�<�TQ������%�x��B���:�.�����g�{�
��#[ŰN���{{D�9�Su�J�ʦ'P��X0�J�I��P_����%�|f���Z���{^d�g �
G�3��n��;̜2̗�Cdz�$���Fh�nI���X��+��޳��ڌ�`��db͚J����,x-ʸ��3� n�Nps��-\Q���������B�/j�����s��6�2�2��8єj� ����$		F����+���1�u�S36�0�������J�*��� d�b��$W�m�o�z�a���\�������k�Wl0�>D4Rl%�{����
�����su�A/%�09�������o<��{_S�>ά��XxZ۽ʰ9' B��~!��Uv̓7~$ʤ=�v3��tﺪ���ې�{n���ml"��Q?f%7�2e��8��2���&L�\�Bbq������ԃ��;v�U�9��χ~/��*���|�n�R�(��&��9G�]h{�ySZ;��^�-d�LJL�H���W\*U
`��}l@��yP�3�\X#���a��ۺ{<8�@RM��<����2X�x+�>nN4��:�����#Z@��G�`�f������D#!@�=SgxU8�|����Oq!̢�ۡIQ�<��?=���onW��BĨ�"���ǐ�ߍg@�me�k���|�R�����_�M��S<O?�3l�D#-�H
�2� k6J��	�J;iH���;[��<o�f�{�i���{�)��W�xH!G{��
|���V2.�M��?�BZU���C
�E��$�Lo������l5o_u�oH)�4�V5��iEQ�d�{�����|sC'v����6뾉��]��{dyH���!�����=����
�$�V�����	�B��f�����K�x%վ����y�õ���V�D����;��EM��+�tk/��w{\�y�c.4�!���� ���up3:������SK���Ӳ����L�U����&�9ŀ���|���.L�����D� ��b��#�*��_~krS�L�ď��h��pWo��ۯˌ�ޱW�8yw���㡤`��`��ŭ\�7ݭ���d���&���*m�L� ��8�~+-�����)�c};�X�\?��v{��#;�n"N,�d��(�������kr���#���b�5��I����s><����夫7޽��&l��;����������ZᗺW��9.o��vq������\�R;`[�ǳ���,�{��?��L���秃���D7�T�]�{�(�9Y#X%�蘻{����7F
b�q��j�N!��9�{kþI!j�a'�̶Z�G^k�I�Q��F<���dDMʇ���9>y�(�Ř�ʃ���ա�s��%`����Z��l�4n�pVdP��= [Fg���}@uI�:3���~J�(�M{Y��PQ������R4���v��!���H�~����&���B�D�	>�>�j��)t�Yl클����{U_X$:�:���J�ŗA!����[?Ы:�ъ�� �1e(���Ó&�﫸��L�����d��%�!����ʆrH�����jVmg^�r@�M����%9u���[9|��I ���()��߄�bv�n�-�-G)p=�����n�z������9՞1�3��?� 5��o�RR��ݿu8������ɡ';�[�Ȫ��P�^�����r�jEz6�zT]�XEf��"�.	�wM�q�"���Z�Μ�^���8�WI�8`�5oz��eh�f���ȣ��~� �茽�H�wv�\z�{u��;������\�H|�ЍD�'�Հ��&������D#�{ԑ�s�Յ��QjO�.H_�(��J�+�~�2B�f�V��f���2@Y�\�M�|�]� �O��<S�&�����z!�"a!��7qenG&Z�%���}�Q�ec��kr�Z����x���	.%e>7��^VZ+2N=+A�S��<��fO����/��n<Ei���6*�.����Z����#��o�����sV��b��9�I,���^�Y�l���4������o�|�z�;Q���ng����痶�zZ:��������)��Y�ť��7�\�Fʏ�W?\\	i�6���K�����?U<���?�zF�/�����6�����jh���K�k���i˽�\:m7o�/�_u0.g<"h��.�sv��N��1�N�>�ɒ�U�w�F�dH~�if��[���M���f���7O �=k<[�ZVV!�М��O��U��o�>r���i�C��i�^�[8~:1h��]N�vh��]�?^�>M#�S~2g�B�ZS�S_�������-}}-U�r�j�!��ky������q�&	���8�W���_��y��c���)/�yz5�H�����D�{a���>*�ԗ��=�˘n!�@1z6xCy���wB�۲����N�v����S��:�F����KO����������iyt`?Vi�V�G,�P1D؟�7�*���ZDDI�	�8�}��}ʁu���F��@��߽�O:h*��Вb&�}�&����g�������fq�Z���&}��PEc�9��u���X�v�S����K�$����P
B7�}��[&�_W4�ֽ��a1[���-E��6�����k�M����1��$i�E츺�:@^��e��Fz�7���gAj��|,�vJ��s�̎R��,YY6��&�&��<�l��X*l��*%с���7�����Gs_�V�1�݇�t� 庴ՙ���9�����gꦏ�?{]� OU��rR�PL&�v�aUt�N>��΅��V����}�kw�%7	���7ݟ����N�7�1%���f;��,v'�$q)���S�A�� �zaW��z�?���.��5P@���)Y��MR�������Դ�6�ч�agP�&�[a��6��s�"�լw4���;���oFv�:�$f*��տSZ|����"��vSgX~���޻�}�gJ.�A/Gm>����Q،�ע���>�s�+^^]��s���.���������=�(}@*i��zX��e ��(ў����6��z�G��ХWN��o���8�ZJ/�W�*�>����ç��+��zN�C(��03�.�Uܬ6���m,dϘ<l�Q�����(54q�E{��G}��㋽�����+�^OM�<�����eþ���`����}�N���u���|{�U��`Σ�vv�����x���~o�)0� {�4�g8���b���h(j�VJծ]��ъ�[�U��E�Y{o��3Z{5�&�h�������y�y�q�^�u����u;q��?-���˕u���{�~�GmL��j�r�#�LT�̆��WETF%�Y���.��k-�m�����;<�X�.�ΣlܣGw�s֑�Ə@��������G�8f�Bt�i%ݟ��I3�WxHŝ߱M��v+O���)Y�[�����W���IΑ�sÄ2�u������V��4�K ��h�O��`��i���N]<!�w���Ы@�H7Є�J:,!p$4(w@i#!��Ѕ��(a�RN	Z~���RoyP\���7
)�+����\���1`�$8�6*�2#�Zb:��I���N��i����U{J�l�LLC��@n�e��@�Z|��\�����}�>N���׾�㱐��oV-�����I��ԗ��j�i��a�[l��ۧ894�t]r>�[U|p�y?|w3�r\����=\��"��@ѣ����`�{#��l瀟R���D�-�p୆�Pm��X���s�� ���MP�~����-eC����d�f��*]���1�(���LA�R���$"����a�ED��[���m�.�9��*���$j	ݘaB$�x��']N�������G�;�3\�d��ʞB�L�d�� �(`8�;,6���i��4���½ꅫ!��C���8�oG�%cω`�_Fl0�D�l�1��w@���^�h�nf�p�g�?xߖ�%[SI��a�kBn#�C��>	���t�Q˳���|����ە�P(a���n5��y�� ���S�������1>X˝�BK��ߟ��.�;��'k���L��+�P�^g�(wɟ.��Dw�p���{�!?$��A���\_
������ѡo��9����C_�MZh1�����P.$_�{�>_�c���B�z�ܨ�y|8w'=�y���=�s�m]��;���O���j�FN�|,��!C%�=��r]0cs��O��Z�����4���y2�{i���)�|�'Lq5ے�=*nq(kb*�'�r�0t*^ǝh��|��q��T&T��x���1O��_���&���!��ޗ\Ϝ��Re��9l&�B4����aLUn�à���ɋ2J�QP]l��ٍ=��|x�q�ԛ���x�iP�3B�u,>��tI���	�x�o����h�xvDiOTr���K�*W�P9�fVBiͳ��������s���/�j�Af���4aKi�����#�$�û�?��=��^�A��x�ؠކ�if;v�1sT�P0c|xh�� �3W0c�o�L�d��^ay�Rd}�4��8���#"e,�C�g�h�tjY�3��u��g�+y��좂U�:���R�mqSwq��EME�"���]�3��U-#_l�m�{���j߯ꕛ��*�Č���ZY��������������?��^���_P��x��=�0�x�Fm����eecӹϋ�?�f�8���P�9�54��PbL�ܙ[�ߥ�Kgw��3VnC��w���W��c�E�O�T���7Df뭔�.Ǫ���w�X�*�+7��P����`�vJ2_`8ѩ�
�\5d`e��ueЖ�:�)��]4�灩i��мp�E�"Fk�AOz�-���u��C����N��r��M4�����y��1���,G�2��M9J�N�uaL��Uؽ�j1�즼z؟#p�q�lJj��DC�X��q-oFMU�����KD����#.@�گ���vo�H�N��Om�6�am �̼r�>c#���ULnK�h�y�� ��*e(�-�)��ѧ��GC�'�vU-���v��ѐ�F����i�β�ى���i��//%�^��xF���Ir�n�{K���)t0+F��J9}lJ��N�өE�#Ͷ����v��4�����̹��l�l�y<=���7�^4s�Ur?g�R�1a�n��
�fA��Ǚ���G,��?K�0�Q!�L�7׌W�p�@�]���ٜ����*uU�.}.DvP��/\sc�Y;MD媓��/DV&[��#�j|Q)kL�����}&^v�`�'&��)(�̚�{XD5n���A�D^�X|��$5�>��ޱeg���b-[�@24Q��5��I��P��0��W��6�iR�.���rB��<?�����w�Q'kr��ß�'U��%���}�����J(Ց��v��� �F��Q����{�ܸ���X�M�p��?7��Ʊ/A�p�]�G��� }��̵���?xj��u�����GP�G�"�xgb�y�&�F��H��T���R0��>�y�t�,'�ʝh$+�/�ו�;1�6ހ�Q�v�_�T��&�A'Rf�O�S��º��/�B���%,AS!"��gQD�Ki
�(���L�6˯��S�	���<��L�~�i��5Ã�^>�] z|6�>����*��������P�_V�����B��\�0$+�F�7�E����Gп�/k��"<i�X6U���~�v��F���_x���%֫�%Ճ���e9<��*��h�/�wy�ʮ5��9�>��>�]�@f`�Y����d�n��#��LI|�^4{��?oܪ��sOl�N���h@�.D�����5dS� 6�a�W�8��9~3�gw�Ҏ/v�y+Ag��F��+6�Z:���R�T�F�@��ǡ�D�!�%�X�)2�����̯ɚ��/O�6L�N�>Q�Jj�Ċ��]�6%���t����{�ф�i�5'����+��
�!�f���W�T}��ۦ�%�T��h�����樅הΨ���PEp�.��-�7Q�����j���G�E%3o_�}h�~�g��%�i�t�1u1K�C�V��O�v̡��rN�����j�%����C߹ A*�pf�#����&^����O��X=�?�[t����c:l��y�g>�����=ۘG�.Z'	E���.���N�_'j��We�����L]1�j$�?��>Sֹ8}�#e�..j��?U��{m�;�(��9�k�(,�B��)��U����0/�ZI���@3�xA�qh�D�k�i��js��=T�aP1m��ޮe}X�A�#ׯh�߮�p���9&l�Ֆ�4=[��Ni�Uyo�MV�&'j��N	���z{���i�JE�A�Ճ�,'�p�����q�M䳀}&�roè�?�}�msW�uZ����qm�N�g=�;T�H]��ܙ.Ob���}�����S�q���E,4` v�|�߲��F�����5�Y�g^}܅W�?���QLoԿ��O���E|��"_���9I( �dJ^�ܗ�&�����B�������T,��w/�@H�iÄ͖��P ���E�b��4���Ɩ��<i}#XDܪ�O&� �J.2�Rb�����Q� ���x���c��o~޲�3�� c��6�A�N��J���cI���*T)�{^j��	 ���ǚ�+�1J~�(o��른l$�����`5ꢊ����ʲ��뽣��Z?�q[¤@�\�1�ݵ�^��K��-n���BG<�D�]߾�V_PK7G�r��f�ȍ�q��!�A���ar����k�H�D��/�����>�H����!O��5�Ё�Hz�m����,R=�xSj�Xme�Xޗ�'��K(]���PF�6bg�����H(e}��i�W`=��tm�)��}��R0���6�QW�B��ɸ�ReZ�w�
�a��ycj��A��B�{�%���R�Kݱ;P�5�YE�7�M��F�@�������%�׍&\O�M[�M2�^��)�S�J��%���0�n[,ҔlHy>�^��N��v��1�l#Ω����Ͽ����<�
�Q�X$7�m�2/�Z�v���Th�lr�h��J��8�� &����>�͖�;9����i�m�����Ž��X_�B�v�|�����Z3o���T�Y����Ņq^��pF�����QN2��HuT#�U�ݮW�'��}{v�-�W��J�5����<���^Ɂ�:�y��ǥT��=��
�8�F��K��.����z��B�����up}	s����I~��^1�)��lTx�'��i�U1Rg��Z��sE�\��T�Tq}�%�%H��ļ��� � �G�`<�[�8]^r��P�_�Z1bb�e�/��) ��[����C%3%�|����vmB����ȿ���Ƒ�ͣx�����o�6�'3;k�������Fj7�7C��(�PuD:��輚��}�f�<��ܪ�����=q��nJ�/��R}���¤ٙ��ɋ�n�qY1W��� �Zu��Gǯ�1�O}$?d�'�7��,�]u޴���뤍fK{X���&�=��ݺY��Ո7y�y��e���R���S�0a=�#�A#i�<��_���	A�,�̡��ХR��i�L�0cR2!�< W����
Ii ��x����1.4-��=�����9�,�T�9%�w���I�'u�\E���p�Q<yjY1ߢ�r�����'/�`U��k������b<�)��� �`h�+��B��:�U�f7*qY����?������V�_���%���!LܫG�����J�!�2}� w
�v]���rT����6�I|W)M�o�]����J��J���~2ћ�ݿIL��u�����ћ��%�ʷ���ez���V��>��]ܠ�v�깾�}Li��D�
*�����Ձ���lc%��mX���OG8���MN,]�T2U�M��L�>V�I=�\�銲F#�ո��ל����ve�ʜٻfS���s��iXx|8!�E�%���MŃ����(Z�*��w�´����;���2^EHދ�6�A)��\=t�S�!V�"5� D'��G�d�B�`v����5�r�y>H$�6w�X���T4��F$�	�Ϗ�V'�)	p�ga��L�Q����y)���#T+ǛC5��{sM�
�qW�LMrSd��!B����j[�r��y�g�J&����q�S�n�d5�LX6c�r����l��~�4��ˍ���>���������%d����$�0�q�Q�9�|��+w�{�Y'ȇ����/�x2K�i�(�`?X��߮ő������ T=��b�ɰ�Xs����$1�ş�\�8��{JIs�x�f���"*��0�!��*�QG�9�8���ǼJP ��1�e]Sb$}��nx�K������f��l�l�l�C6H֋Ǐ
�`X��^�2C�750� �Q	�H��`|��qN_��N�h�����4c�ex�-s�k�8���~�dz̕�O3c����O���>WI��ko� �?͠Z�t{sP�� &�0{�RI�i1�-MR�2$�6j>m֒�-i�F[DBݿ���M�g�M	��8$n_���Vy�'b���b<O96={Dx�y�ʍ�vM�����U K��?-�)�X�u�����d�ɣJȘh����O�mUn����;S���t���&zm^�g3߼y�����f�S���y���<v:R���P���Zr��+��3'�帊̸�.K��x�g:ƑM��<q�w�Cs�C�YG��9��Kq��~2X�²�Z����|�|p^g�З� ������"N�q�!�/� R)���#�p�!��H}��*<��9�I鴾U�3V�6���P�ݕ�:H�ŉ�ô���;�c��Y�	4���_�x�a8c�g�&���x!�u��u�βi���!�Nm����V��Â��|P
J��fX.`���Sm{�=�Hy_�.@r!� ���ʜ��׶{Q��R7V��6;L��ħ��s�e���݃S�΂�����F���\��I��^TB�����йoJ���>տ�|x��vL��~�����v��J�EƔ](3J�z���~����&R(竼}�C��E�z��^��(2v���u����T���G���Y��L�{���Kd���!s|�_�/ �|$d�H��>M�
�d-��&�q�
׃s��t?��]��׊/nʮ�ǐ1m��1���#œ��w��k�'m�)��]<�����5@/���\�M�#�A�D����j9*�g�uW�V��Ѻ>8͖�+i�,U9
pS�3�R4٘t�V�6�
l��_�����%Ge�3��Z����B��t:�4�]��ʍ	=�r���~���QZ�k�k�]����Z4n�Om�N��(Y����@�Ѿ�'ぺ�&^y��)=o�'p
�:���$�w��՛ˬ� ̍(ўU�BAӏg�	�|kމ��H�,c��C )T�y�N����\�Cʿ=+������6�55��)t�� _�a N��|D�2Ÿ�8�lnJ����P�s:*~%`JRւ{F-uz���cn������i~��k9V�#���M��B�W���Κ0�њx��;$�J�z�I�����9��=�%����+��bT^���e:�|�����/ISXM�ڒ	��2��d�;O�2��G ߠ�B-3'kuo�!���b�5����r;��`���Q��L]���~����۝�|UQ�Mȵ0��LU�U�f|�mV�W��!}C�D8�[S]���ӄ�%26Kٹ�Fj.s�=����3�y
�����Qσ�w)P��06��M�]����=���WN9aȽ������ꫜl�ؔE2��=i�B�^i[wԔ�y���@y��݊�{k��?^�
�i�Z���K��p�k+�41��=����G�0Sc��A��8�d/>?$2�<�i��|���l8Kni��L�W��Rm��H��qM�^R2b/<W�>Y���F��v#R!)���n ���<�f�x}j ;�b=c�ޚ����8&���"�:}�2U�i92z����y�ԏo�t�~�}���A�%���Šx�94c�"wU��Bl�/�|��f[(��@¼L`�lL���MM(.G��9�����R���:�	��$XR9�zs@&1J�m�)����,��*!	��Rj��9=<0�$:��GM\�.[�Ϲj�^�����͈ȋ:���W�;:ˡ�J�'J�-��X֩ x��r����.��p�C5ͦl7׽�]�w��вDۓBF�2:8����f7:�\�_�sE3����O��R�l��c�[�wuh_������݅���r��K:�uU�7�v�k�N��Ȑ�u+��
Npw�X��������T���^X?���z}��˝J����n
��D�6�ֶ���ҫ�ٞR���h�+R�#�����P�.��~|8��s�j�&�^[�j��7Kr����u}n߂ز�X��p3�x-�6���ul�L�6�x02d�Y&� ��շ��Y~�ѓ"�<�?IA��	S(��#�<�U]l�$�~�↖���;f.��T�m/t�\�ϏR�	M��5R޶��|a�ag�?z�"p=�t� ��$�~��Z�����v�+���ۦ��j�F�O=e���x�BQ\^��g�#�_�z�U>rK���F�"�l2����M���J�v'��+(�ˊ���Ci�A3 ����v�����߼��"���L1�~�׀�È���6�0��'i����uj�ޱ�
���(W��0F5��kds}����Z�1��^�ee2�Z�W�.�u�Sn�e�u������e�N�|�}�u�UZ�|��̀�4���u���RXv�)���ܸ-���#�����%�&+c���R-شL�@g%�&o�M�Aݳ�j�&>���b��
����!yM�'��y�8�P��.�767�!�G���on��e�듭�ڎ����!A,�B�"SA0:BU5��S���qչջ�5.��OYx�3����ٺY��̲�~����#�r�ity'��D7���ׇu3���=��W��<N\�G���Wʩ����/�������|wL�v>W.R���F%�h)~���{L��x�Ζ?2��6$^���t&��yc�!�����������c2���<�5����3\s7ӏ�jR���WO��	� �r�A\Dԛ )<jY/B�.��^����f�����dr1��iC�RB|�$�|����9uR�f����f��L�>/�ysu�x"��|}V) �Q��c�>��v�Z��m}e�ȥ0�@����$`F.�l���o�/OND�<��{������Vx��,4}-P��
&�ȸ��六����]Le0u��`�����}���{�t�Nu  �C뉲�<@R���,*އ��Ԫ��;7������+�n�����x@s���C�\�W�9�)?HX�g�2S�%E����U1��Z��u6��ꋩ�/��P������@�B�V�6�Q��CSJ�7�L���9���"�3�}[��W�8cѷ�>_h`5<���!O˂l��54�9��p�ދJ�3E7�m/�CX���]���ٕ� ��,W$��'V�����@�{��ݠ�o�.����eŪ|���e��l�H�i\�N�]�Ѭ�2r�0��]��Fa�����	ɋI�=�)�3�:ܶ��%�2⪏j�?n���}vs����XY�#�^���O������Up����y��o/�;�I��Д&`����Sl	���|�ӕ$T�Ad�,	��rK=I��C�`ڈ}T$��_�b!]�@��)�T�������%���MXi#b3D�u�i��몎���(�YAi^14��"m7C{9�gq�@j7C���&�å��X��TaK�⚚��>$S��t�[���d,|��f�`��A�toiL �>PEx�8~ȭ'Y�܅��X���j9@ݞ���?�|�'��1���y���F�|�<"s��2V�o�}���-��W��
���E�	�=�d�c�-�K���EA��&H����4��w�9/
�ˍ7Ҥ��Qh���W!�'|C�ή\ʏ�����WF�"�Џ�ƿ]u���T�R2r��`��3q�	�x�M=���;�����6�ZK��X�X˾�Gc%�,g(�LEV���M�����a�0(6Q����K����Y"|�iZ�}�R�|��`��rf��Wn*�v�8)��D�N9^Һ���>&ZV�����?�W������Ց�ZVCҵ�,��f"
�/r���oo�ל��
c��S�k����f�co�c��b��(���4��"�r d�+�P�j8�`(���g�D8�r�BR�Bi��=	���<_Q[Q_,��hF�R��^Sw�+�#�����H@?<e2@2�x�#?�Q��#��l㍪Ƀ�Ɗ�~���6��L�������9��=�7��6H� "��8V�>~�ԝ��Z�r���?�LS�c"��,#����Kl�e'����ؾz�$��\-�r5��I
a՞�|(|�"˓W��w �M�:y8�OT�M�P��o���=�;?�-�::�x]��P֯�YM�9͌�^XC� �F�HEħ��-�M@K��o�)�����u�p���v9Y+��ԓx�b~�E�E�WB7�)��iJo�O������Z3��2�}"�Ld��j��~�=��k�tZy竐���x���eێ;i��I3�~���o��Ia*�·@�R�"�������x:�;O�C�n��]XG(����B���pj3F��=�a>P�^n��p�pF}���4A�� _)�.��S(_D�cyߐ*Q�$�/�W}J�,�a;�����3����%9�Q�y��LXkh�p
���o��|>��]�H������a�������P/���C�Ѹ@մ�޾�8���NG�[O�u�p�k��ĭ�友
�� ���^�x�"k���g�T����R>$�2��|�G=P�h����^=_��ǥ��;�Z�g�q24jS�����:Dһ����!�_-?&+X��V�J�����_Ц����6r� �p=�cL�����y�ǃ�x��Bޱ�o9m�oX�\���3��Qh�,��/��bb�� �
�Ȃ\�Pu���;������Q�p֋L;�"a���*��]�3$�s�rş=��]ځ`끆)�3}gKh[c���[��_��\��N9^_v������?��E�w���Y܋����}<�ϻ߃40~3yO��lꄵ�?��.z�'L�"̯��^�:}��c�	���6"�#& �=X��D�#vR�2�K��Wy�R�J�%�ׇ>T(d7d�(a	
'���(�6H'tm��#�	v�"$�#K;W���X�`N��]n{�a�6��>4G�]k� �O�6@�VRG���$��~���>_�}i��}�B��G'�U�$y:*�'�����~����cņ{�B.��&��*� �m��*uI\�z��,U\�]�]͊���`�}<p©�Pa2�!���y��f�UrM�Pl�!Pw*��%�1'g���������L�ꓠv,Z^�oi|���<z{�n�B�������������#U���*�"�\&y�	�go�P쑌�m�輻 �H��_|�b�*2 v0�'J6��ߠmrB�i�;,!/��g��>]���"�xb�4q�(O�@9��R�4D������.j-Z����%pȉ^�eNd�L��g�T�=�@�F@��κň�b,Ĳ��p� 
�B��b�'��	�����oe�kS-���#{�ZKwN�M����]WT�f�@]dj�#a�5�����ko��wg�@�h��r���ꪝ���	OWJ�v�V���AZ۲x��.��C�t.
�L�S��{����>�ҫ�}�M�i�u%���f��~��O%�߯g�����c=o�7��;���:1� T�ȳ�h�O���1ԣ�7Y�����<�y�=����&oz�(���:����h84`%���ɚP�
�&�D��u�}_�;���c���������+x1��NƞH��D�R<��<7wO�����Ӝw��p9��4WBW��ؐ��W��r�V����>^�.�b	Ơe������k���w\��
�bS�0\�q�ϻ����O��p�b��8ُ����{DiK����H�Wh�ˑ�S<�6��r�q��(>�v����*	Zq��x�.�ɉ���'ӹw�h5�tGp=^e�<�'�Σ��y+����$-���0��~�9=�NdXBЗ��[i��8��8M�E��de�	wO���=��jP�I� �9�����cKS�OT�go��_A�ɓMrs�R��ÞU��9X�=���n-����I���@�Cg��H�4
�����!5 ���j�����=�d��v�˂�>��q����Ai�N�?�o�}�]�/Z�ݞr�B�F�� �Í�-����H��V�����i��'Hd~3h-�����C"��@?(�i:^���=%��Ф�����W���B�I�è����R��KM <�򅢛��#A�P���5�1"}:Hr�{(X����oǠ��~�i�%��9�(��y��'��續�Y�U���ն'R���<W!��3J�_l��j:��c�o��U���v3dO���.���BC;BB��M�~%��^��nlk�=@�d���F��nO�l��.Vaz� ���X��w������b���2v��%b�8}�"p@��}OM;�����Ȑ��w�`��?h�d"p���G-��(r�T ���,��<v'*�h�a�)���s���S9�YPeQ�x���O!�TU(��YmsS���
+�p��H�,p��ȳO�E�[�HM����?�Mmx[�p��9����X���=�Ѷ/j�49�O���w��#���ۓ�:M��������p����)]��^� ��g��z��v�Q�@4����g��2�2�6��Ҋ�\�!��LL����� ^nO+�Pԫ�IG��L˱�kq�ی�������u����I��B/���QV���{����mibX�e�m@��m		���R����|%LP��;E:���K1�{�Hk5q���+���s���r�jbS9xm��=&�m7�����	�S���2�t��"W��d�W� B?B����.8�9����{�����4���J: x�� ��iY{1��F���Rd�@��@�"�T#\�z�)8A!���@�#2~W��aD��������^\p��;Դ��om�@f7�*=�:�&��f��o��m��b�������G�';�z9�p�wBU�U����w�e����Jp�'�޻�g&xR�K{��
#��h��
�����Xvj�*nF���2��%5�g�,�Yd��7Y�G@�' sD�T]ȫ@�AKlՒ�����1��+db��)�X���D`blM ���P�@�`9/���:��(Ǚ"�?����$D��[��As�,�q?6��
�eӯ������n�[��M�{��tE�
�ӝ���?6��u+����x2o��,@P��p��=�͞gm>��:i"�z2�aU�x�"dT�=�a��e��Ř�*�z�SC�Z�N˭.�� �91����ZuЄ�'%��/�q@��+�ĵH,LH]���wK[`����ͯMh��P�é�g6:�3V��,�M�MN}�	I�A�w`�m.�l�1
0`e������'�� M�A�+��oU?/>�i�ND8�<����Vq��Jr۫i#�����L�1r���������//��<Ï��zU���n�{�nm<�K��"5ؽ���Q�U�9�5E��N���JUt����.5��p����a����@��hN�5�ˮ���b�R�����R 	k�7O��,,w	�t|TA?L��RxM֔�Z��_o9/���'�U��ϴ���`��L�vH5��m0$��zr��e*n��H�(\k�˽l��0��i9�7dLf؎�M=�dK�S��X4f��� ��P�qye����vH���S��4oD��}�~�ѓ�d�3?O( R�(��p���?��mۡ���DlZ|���3��A��S��O�3c##�0�.C���2�H�,ajps׷UϿ=�w�	�c��hжzr/Vh�2�<������B��yA�#�=Z�ö5�y���rT��9�X�m���Ϗ�n�q�uH�᠔FW��Ϳv���AR���pz������ɒ:�' ��EGIh6��`��gvؤ�������=�>��=,�q��o��O2E�D���(�w���G��a]J9�?�J*iL��j,,m�u(U��`k�A?G��'�s�Ӵ�+^�'�<�-ݨ1RORwR_/~�T�z�����)k�-K5��-� ��
�
�a���Y�V�%��v��A)FU�<R�u1�j��)ȨG�&de�48%��iU����>N��j:����HY"j�ѽ�S��p���oq �Dq�Q*��6��liW���Y����/�����������-����m�u�.��/?tD��[��4<��vv�e���gu?=� ����L��W��O�į�Y�"����8�W��;,�%�+ޟ7ܽ�u3�L�0������)r!�¸���5���Q�����W�26���w�S�����i�`�)n�!��|W�T����9���s��u��e"�P����"�����=�1ƀ�"9� �g؄�1	��}��꾟�/F])[���PE7�C �f��tI�AM�����)\ӝi�R�lV�ӝm�;��zSQQyok����.����d��S��N�W��S5��?E��5������Pp��B��O�PZ�-�}p���o[D�|�݇���c�8ri>�@�d�.5��������i�h~�dy���i+���S�2���� Oj��g�%�A�l����[V� M;��h�e�J߅�wʀ���/�ŇZ�|]�q� � �_�=��۩��)ؔ�<�B���¸��
���u%�����F�o9���blˏ�XyA48�$�mִ-��(��ioL��MT�G�,��~/��UX����Xt��f-��H����[#�K1|'���	JU/r{'�o��m� ��#""4��e��s_�޾=�����Υ�|A#1�B���82��W�.��~��~���m� �T9�� E'��9����*8�$x��U�{���Ҵ�L@��Rʼ&U�T��K��֑��	38�[��"7o���Q߿������`S��TJ]���c�d~����o���F&K\6��.`U���]7���"-��N�D����!�$`=�Lw���de*��ݦ}sW��f��7-eV��?�8�o�8�?!^�����H�L�[U[������s��r��z��8r����N~�@Z�e����Z�)�X�?hoV!{Q���HN|>�詖W8�W@ 9���К�l�QR�'Mr>%����\D��#$�����3�b}���s��~�_�!�<�Τz����������âɃ.m�p��<�;XZa���.��X�Jh4�u���l��9(���Y�;*��b(Я#<������${�4�>k�I�X�>�~��):��9r,�ɇ[s}]�wTo8޾~�t۠��m���s�K��]*�Eۙ
ӷ#9�_�(���������#�B��M�_�M�}M�IK
��r��*UN�7��*yOZ����#�cr��6H�dp6C�*)&s��f�?�u� �){���A���m��q���Z{{�)?� ySJ1m�O�6�Ȼ0���e��i���Ln7��k;��J���-��yA,^�-L8��1\p��N��$ȭ 	���[J�
�y|���iL\�0��l-��;�p�L\}�|S'Ȅ�z[�~6W��i��N�^d(_��_|�oq������\���a����&sF�Ph�j
�fN|s�l��r�,U�U���<��L�N���L�n�M���Y%JH+�s��½q����V��_+���X��ƫp==�6y�c��,jt�TA%~M���Pr/̃n�m~�u����B3�N�A������o�h&n�8}y��r����O���?#��ww{��3�r�v��_�}����H]�� b��<�8.��nԥ4�'�������D���չ�E����_���~|�m�t�
O������]|��{����j�9��]�6��� ��(�T{n ��AD�{�R4Z:�����9־��;j��-�9��&�7�����0���%EKS��DT���wJ����c��9�N�_����§3�l�ۈ�����J۹lL������(�����4�-��Q�#�#u�����#t{��"����������_�m��r�eO��"���?��Ö���o�vQC���)Z6**���@fZ��ܷ�֓@(K^�c�3�u��H8KP�z�X
�JL���&W�4Q�R�1��{��x ����m]�ێ�`�n�0���I�N��ꨅ�ۮ�2(lg���~(&�	�Is�F���";U��;V����Y_چ�I���ۘ.�u��ݛ�/�j����4������2{#Y���A��/'�)>�~�Nҿ+��D�|��W���r��Ո�k\�%��i��n+~�A�ġx�HQ�,18�:%H�A
 ���eq0~/3�p���gB�6R��fMv5ݺI�аi"���(2��@����h����9ʣcT��Z�R����⥩�yez��w�ő�u��Ɨk%�>�ʧ`j���VdAx��ji|����Uc�~K[�� ���
���Ɯ�$�$��.׫��_-_�L���h�����|b-��y������Ҷ���[��a�8SsL����rH�7g�� ֭.g"=Y�-k�uJCX�*B��� ����St��`d�vݦ�utp���LV^��|��U�G�2,0�﷬/�l����jLlH%^� �͞��T[��طL^x���l&�Kи��q��R��dt�hׁ��}�]� ^�Ҿ�����޽�:�7�w�+�؆:����̌|��D�������R%�{f5����X2���PJl��  ��C�,�,N�<�d�
�I��~C3>yԕ���]@V!�dm�@x�Z�t^'l�7��
d��tl���}�9�q ���&PU�lV'4&�g�`��K�^t"�/�'�_�E1���-�d�}��hw�PȤ��S� ������4��c�iq	/M}B'���9�a��Tb|w�bC�]�)ZoL�m�������yi*?���n�i��o���+{a¬5��6���i��B8�k1�I�'��F^a�LS�q���!m�[)8�wYk{�AJD�J�Lm�+�pmL���X������Z�5O�������rq㰦��ܛ�7��#���cGr�f0)�R����(���_��7[}L���^�vq��nm�����?^�}d��>W�%�܌���O�j��V�	�<��H8&p��w�ۏg�<ZU]O7��vE��x�KI�PwFjj�g>j�Q�?�C�x+�6�瞪�b��Pp�vhY�w��K��W]��
�%�������M���w퇂��a�[a	��b~Zz��۝�A	�珇'��Ŗ��jl{��z0v�SNB��^].�2J�-��{�8�;T���B��Т;�m�풷����M�>��᷻-�fc�
orP=����R�j��Ŷ�����?C��+���y�v�Q� �U��O�M�rAhǐEQ9�",&�Д<Q���E䧥��K �/�F���0qK���c�p[�Ƭ�w�E�Oioe�G�2C7���4H	*J!ҝ�t!��t�� C]R�ҍt7��w���9�{�=��5�u_�������*�j�ƌazCz��}����J"^.ҿ@-�뙋�GM[�6�H�osۛ6��9����"jf,1r8����ƅ够%�ܒ�7��`ď_��Bp�嶤�n�d�&�r���$a���O�n�_���3~]6���xfQyCȓ���<���x�X��)�0��]d���y���9����bcbNb����Ƿ�����4�[�9,�ъl�u�+f��
T���bM� ���:N��~�y�f �J����YCCC%g�}�/���\j�5�}MH�b�>�ί���ը�+*^��9)&4��
B�-���O���]4@�G�O݇$8�D�9@�BD_^_|������y:��gѷ\��տ �ՙ�|?�x��dcc���lA�$񲤇�#�7���a�Y_Rq$s�g�)��ڴ�F�d80Jyx 

�M�`�5����<���L��Q��:�{�LkAdH�d�Ŏ�}^�u|�\�r��d�������$�Uɰ�{���(%��a���o߱)�֑�R�oYM��0�C��kќw�(�6�~X�Y��v�Q��ӕ�N,�v��צw��H"w�K�6}�r���b4Û�`+��\Yb��;�>s�>������[�=��ڤ�(Y��� �b� ���Y���N�5�����v�Ւ
ė�_h0�S�<�19�К0Od:�� Rψ{���q��,�S�;��Jg���%(Խ�L���nu�Xg@dڴ;Li	5� ���'r���V�%{]m�O��T9�G%�A�5�@ahB���Wi�C�n�(�7��'�W�����k!�}�kyoC�wEQt��� ���)u?\���d�T�x,���`m�@���$A2|4����{��M�jO����?Hȕ�%�031�:���+��N��`h�v]}�_"�!H���1> �hR��������/v���~'K;��:U��=�J��[�fOs�;�Q�GL�!���۫@�Y���NDŗ����I����̪�Q�r&�x,N��V;[���|�Hx�}{>u�Tߊ��=&sQ��;����H���z5�+<b�Q��5b��-Wd]��=����O����?`O�^�a� �/�^�E���RGj0�%��\�z���d���<�����:����3p=v{
A}�:83"�v�O
�G�ϛ�jp���e�᫙a����%��7@?�8�~�w������3�������Kg�p�d�p�n{��.L\)Up�F��*�a5Rx��	�+�^���׼#��i�Q꯷� W�k���Z�:�JאF�‽ɑ�#�kd��:6���ҹi+�:8e0�zO�t�e-���1�P�^�OnL�w��k��#���.��۵p�rh��F���.�a�+����芘b�`:8�d�Ϣ�ԭ,��O�U����$��-��4����N�%}���0��u����Ռ�B�e�n7��w�%�ٓ���ii�7w�w��%��e32�j4���T<��k�`�7EkA��JW�I�:&~}bs�D�O`�1���'�����*,��>`�G)Q�]Զ�d��W�Ts\fuj`[T��(�`���9�c镇��ԑ���3P�ǀ-[%�e����&9����|Z�1�1/Fr��jذ�&p��t ���Jr@2� ��y�@z5� ����v ������t�eVx���q�X�N��Q��,�1�i��n&�C�3/g���Þ7��Y�J�����z'o��0p�o0�6��J���D=?8�b�H�w�� `{��1�vk�@\|6��r�f��tHrQ�LG0l��l�DX���HB@��L��i\��YW��&�����	y.3�D�u{s\ޏ��d8	�z^���e�j�a�\b����"��N`�w�ϧSzLuW��O�� g��w
�--�&�l�6ʙ�M��5U�5���c]�(��m������%Cb����+'i�6Y�-��m��l�+����$� x+��_�ͺ©��~�����<��:0<{q�"R�n�����<���nc8���x���r���0*K�NE���K;&f6�}�`�t[ۊu� ���MNR��7!�:���]~��`�����GN��X���:W~v!sIȓ��v���P�)��U�Y=�:�|�x��WH�
�p�ҚD��������bHh���U�\���k
��7�C�}�ú{�v��BnOD<��0�F�� l�3W�a��  fn�{���"�.�j9�?%�e!D��� ���B��l�(ZE>Ha&R���T����H �ͳ����Vl.86�W���v���6�q=f�7J�vR�G/ �Y�j��@�H��M��0h�H��DG�A�SL8�L�?5N��R�)Zm.��Q\=(~���6��I6 "��E�����2`d��)A�������!�%N=�>,�f� ��n;����~��ҏ	���w�k_��4��vb�7�~\�`4�ޞ;��]�YO�O��]e$��׍��h�n(�eZ�k�Ѳ�s[p�FN��M,xn�Lh��n(�L���l�&8���p-�A\�v�_��)���C���҃Q�6r��E X6C~n�Ǔ0  ��Mɍ|&I��h_���5#���[��Ȓ� �5H��G3���,�e+"Ȥ�GHyyOV{��b�<c5�2����@�äQT%#E�6�����·�O�ah�6�~�i�<��m?rW���l��J���#���1��
����U8k�i����P"�u���u�H-��ǛVtb}�j��Z��~�v�?�h9'���z��1��g+;k�S?��gf�z�	 ����\âf����U��~<�K��:�׬kO��ZO�l���y�Ϯt�D�w.Z�0ύ<��͍䤫�"�������e��f̈[E���lǔ�d���$;�^`��2+�m�6%	S�[[q9�}%��#�G�t�B��h�#��Ѵ*B�]Vt�wph[x^h�&?�}������U��Y�>�=���N�0y�������؇T��"d���`�02?�p�����k�e��o��V#�g�+�nlJ��]`����Fx��;�62(I{Q��sV3�:�i�����!c�0��_S�x���wA�-�wLߛn��Jd��K��M��U8�aB�S_�2��IbHWc���Y�ylKXM}�`Zf�_��0­�I�+��W 	��b��G{ti"��X���_+�(��{��1j^x�M�*�+_�Oo�ſ�J��a�e�e�����6��<Jfɦ'��{ �7�`�׺�WI۔��#�a�F*�s��xm��[$b���X�[��L(m�ʲy���\[lηV�=O[�ޝ勻,@A�"�;Sȕ�[�%���<���?�$͕�� ;�����qQ�YiEmA�P�������G�^B�n�w=�R�ɸ����%x8qK�1jSʵOp�� "1���q�՞-]ӄ/C[��+⑵���<J�-����g�d{F~ߨ\0�"�f/Θ}@��'�̮}���FҘ,뫩[>���n�S�si��FtfD��_%,�mb�ß��;9�d������8�����0���yf�JB�h�ޅiΤG��@,����L�j���|W6���f,���_�����K>��܄��F�kz�]�fާ5I$�W>�p
�kr�%�Ӗ��]�X�g}���lK��.�����\��F�RTV��4�"�;Ԭ��^Z]��$,P���t`��-���D���M7��	d3�I��o"u� �1�g���U_}L{�`$g�t ������F`�;��/2ޓ��g.������C_�ʣ �q�/}�Q��Uzy~�������L�x���*��#��D�����AW<����32�y�"�-����$^��uB�!u���:n�5k{z�/h�D>] Lڕ+��΀F�%�������H2��1�FK���\_r�f��4�H�����f�N`�i��n�ot�j��z+A- �55�#
�G�7Θ��\�JW�D/W޹k��8����蔛.e#�N�ϴ��vc�mΡ%Tf"q@�{�����We9z�����*�d2$����)vZc0Vn��E�vg� Ԣ��l�9������k�0sbc�&�
iQ��I�ʔ�'��Ô���;���FG�� Ɩ�ԃy'B�y��MǤ���J�/#�Ӡ;ٖ6��fְ䅼DÝ'~�0��1ǩ�-!�OtP����݆]���{Gf��F��Z���;/��_q7��k9_�[:.-�v�Ř ���<lB*�<ݠuG�r��,&��i�쪴��p�����}i��,أ8	�F"��n�p'������������4�@.�Q��C�-7'�Q����_���-@�y|-��dΌ�@Oȹv��ǺU��[�U��NԎ)r7�w�}�J{�<��t>��9ia �o����mY2<����
=�Wm����Ck$\i���������Y9Z�o<t�;Z��M;]�5�f�Ͼ� \�a�>	��lkX�>e%��=y�3��K�o!��]2ޘKÖ?oV���3�[:+�N좤��{#��ź���J��*L��ݜk Y���f�	�z1�_�+�2t�=D;�|P�,g7gQ2��P�]:h
����	4ML�9.��X��:�n�6j�!�-�����L|M`|n1vqA+�37�f��Z�M�0�0I����z���W��ȭ����7_t��ά����a莕��Ӹ,=��E�I�� E�cj�Nc,� �pYҖ=�N��3�6;HU���]�f��"'k�{>!ˬ���+�w�����:�'��9���]�}~J� n�uD����� b�WNa���FGgZ�S7�{GX;��Q^���p�$�+��e���1�$�򓐨ө�6�A[LU1�KD���=�س����'mElc�pN�nH�R�r�~~3���o&�p���B�z腪b ��u�e�����p^|��軥*R����_Z,x1+t���)����!K�64{_�VcQY��p*x�F@��l�2ڐ(�Gǌ�e�5���V��;������'��Λb| ���K���>l"v�����,Tx͖�vrAe�6ڳ�!K�[5��嶢d��ic�f
���Mg�~�ୂ\	\D�_ڠ���NT��?+�d�3D��S,���z|G�B�g�9�S���6����k浘Y�~?a��A��??�B�I�w������T��zg���q*��XX_�M��Vc�ԚZ�`S��z��aؾ�y,υ����I.q�2��\�����F��V�����ϲ����x������y�nJH��g֖'f���2��;�gc$�>sk�p���O�"�_�д̋�����4]�6�y����9�Em�Gɩ�;��!������A:���f�$('t~�N�V]jc�b�9p]�r-k<2���ޛ��(֫��+Yѽ>�6��Oul`�[ ɪ8�h��E0���������'p�����;xF�Y��O�X�*x#�\�qƒ���z_�����/�Hk�t��t����ղ?zdmf7j?A��mǣ���=��E�^H #��k���k*q	�?@�S�����ɤ6/Vˡ+cQ/��B�G�����qO���h�Ũ�&��C9x������?���(�yS���WM���Α&^�ֳMi֋�֟*��>�}h��aq��1�&�;Zyb!����M��Rq�ij����� �"��uδ!V�z�A�IU\/�����������ҁ.S-r�Su�u����ˇ��T���.�]7�~w`Ӻ���p���f`Q�ۉ�?�/a?�[&Te���_=�p:$�-�| ������u�U�K�T����0��4�¶�rc7��#�5KU����'��5�@���{�
��gb�{�}6�mIF�;�f{�f��|N�Ճ�s�
(7S�BBh	7�5vD̮�b8�m�o�/���z�SF��V �$Z�2Aţ��uVo���8>sa���#��J�|�ܥ������>�ڑթ�#�ԋ���~�էSB~�La�Q���eL��E5�Ϩ��[����D�����J�'sF������=�`��s{���Y׷���m[����n�&�V��J,U���w�ݦ+�s�ra����E����R	kd�d��n3|��>^�]T�5��]���p5��s=�����P�|���]��A��)��FB��|h���Z�� "W��Q��1��2$f�٠��\���"b��
�^���i���0s��� ���rQ��z�.�ri�|��bָ5�ޘ�1��0O�|p10��>_����B�
:$dZވ��Ż'zf$�	�5�o�fz=1C�`7'G��q
�����Ι��[�_�(����t�J?fVpA)�����o�m�޾�4���W�1�n�ІFn��*tK��n���������B9� ��J�H^golN#��G���F�N"�PAX﻿./��Qw�`}�jxӛ�I3+�L��5-�?�L&Z\����J��I�2EZz_�䢙pk<j"SflK}(%����|i��z���i����3���TS�?�$S�3Qg��=x� �e�U��_k�Z��S����MX	�bZ՞�����_�Y�\i��7��_���o�Y�\�X���0PI��O�:�'�3��X[�Yq�fmH���/[X�	�Jsssw▆���ywBc��1�%�$鳍Y�]4*oДWtU	j�F���gF�
z��Z��]g�x��F}6����p��TH�ue'�_K7M��&#Q��a��.���d�Ԛ�,}M]��m� wz����Ə�u��ӫ���Ϡ*��%�=���RT�Z����న�+#���1}��]m�#��`ӗ���W����L���!�=#�
����/��r�.bIWpQn� +HKMMM6Ff��@]0��9��γ��Î��Q#Q�^WlV��(�)B��I
���ޖj=k�r>J��C݆%i~����A(8�ǍFّ3��e�P�	+$�x0-	Ɵ�&qz`���� >az��EW7���r�_56�V�7/�}@-�v�ޝK���8M�Eо�)V��Ry���vn$g@��#Ε�'ͣGM��%)%)�p�3GcL%!�Xz@��Ii�Ksm�
���4:�$�ߐ=ԙ�S�	��C����9�̮�9-S�-�M}��%/����+�>+������G	�Fd��>{<�H�F�ͣ����
`�����Uֱԏ����OL���[�Sn6�Գ�cEMG�{E����Ê5��8��8�Ҹ�����5?�E�Α��ԈL�L����Iu� ^�1'F	��|9A�#|�ؘY8"=EO��lw��TwW�=�2R+��&�&cU���
���l��
���;[����O��6���n����.�:1�*G�u��������D���+�� C�A�RM���
��} G_�?{S;��BA���<&FA��&�4a��B�H[WO�)#�
 z��rM�v2��1ϪI�`�$㉵��%{?���9�ԏSl���wu��/�I˷��3�����'l��01��P�'v���G���<�u��6_VF0-�d+>��mN�7�����/,�:ݥ�P��u�(�b���"�z��N��*�������Gb:Lu

�r�B�٢���IP�y�Ϊ�����@Q��0>VL#p��e+~_��6\{m��U�0��'�	e:��*x��'Y��/퉍����i\Rq(a��� ����,:<�1١�$���BV##�Fg�T��8�Y �[U.�qUb2�s��w��o��$�$~���M��E���c������^&*	��~h���;�~`0!��ᬤh�?|��+��k4�D�>���$�$ꪥ���L�k���7�_�M3�B�֠��������Y%5 �Tp��8R9�ʚ��K+��b�����ۀN�7������1��0}vI����`��:7�5�2�.����wO#/����k��Dc�#ޣ	��v)��~��~�W<L�6�F�v�����bަV#�λ��$�_5犯��m�c[#C�϶�I�;���ng���qqep%psAlǅ~
�9]I�U,����y�x�I�?��������q
����:��<�R{�FJ�+��$蜱�S�����_3�b]~f��G�foR�|��Vî�Q�?ejU >����Z2��RJ��\�,������<���Fwf���%���H�F�ܷ�6&e/;�+Ρ|+��"&ܺ�F]�d�C+�V�$�ڗ(�����tQ��^�,�����ЙL ����]Q�E�ĨaZg����R̒�
��������V�Z�)a�J��7螉�T=��$rg�j']����R��~���'fh�0B��5�eٴ&�?^����kdF���f�h�� ^tU�$8�,v�f�B�*Us��"ގt|}z�HR�5llWc
*-�QM<�����2��Y���cm��'���YZ�ܙ1���CC?,��76�K��p/؇�n�oC�M/�PV�4������^�힤s��G}:C��1�}-������G$1��
hMZ���U�}U�F����� {VV5`���c-<Wk9�~�B׹S�u4#EN���� �$��?�k���+R]��C	�.����24��*�=?hFK�a��MnR���悌��o�B����`��O0N|/�ތ����N�	�I?D�>[r��a���]�ͪНF���y�Ĥ�2	/*r�eQq����[�lY�nXp_E�T���Y��?G�lʚ.>�=�PJ�� ^�:繙�p1�!���
gç@��8	 n���jK��c�=5s��(�[�b�i�%b%~��$�4�$�_����O��u�?_ɉ���Yd�jl�� ��O�����1���9W�r�Z
��E��y��0��Q��)�F����/�ȱ��\i�A�$e�F0�_xGe��*^P�q�|�?��6<R�ς%z��n��
]�N,³�Y��l�D-|&UvbIwQ�)�.��H9��z�F5�zpR���|�̻Ɨ��w�F~�~k=��k��.��}j۞h���� ��)#��@t2!�ڀ[���u�U��$���A�]���4ge,CO��W$�bAt}�{!Jˋ�@v��B����~	��p��#���ł
N�ŗ�\����"v��;�E��i����zʰ�������p4g�za��3��+�g���S7��d��N��{������|}��զN�
�_��-kYLB`G�q'�4vԴ���~����F O��ޢ;#�¿�rW9�,lờ/~[(�ZkZ��sw?��lp\h�g��x�^�q����߲8Ez�2q�Z��!6&f���u��g��%rkl֏j�1�R�M��I�������0�̃/D�;�;O$��I����uV�ߞ��(�,�Wfz��dn'Al'�9P���_��SK�(�Z�55�/�K�r�=����*��(\�%�(,-:5�^���KX*�I�~�O�����Ύ�tT���(>$1����4�6������V)�7�7a0��<|�/�.��	��4{��w7�(OǕ�o����%������~+rN:��Ꮨ��2�c$������d���~}�Rl��n+��vy�?Oܧ��2<�S7^�T<r�������uL�	���p�"��;ϯ�c���f���?@��=k�ݟ��t�e��.�Ӿw�kI�J�IY�y��T��U+��$A�ٕ��n+�}Q�o(��3f>�N�e�<IQ�*L�u^C�=]6o����5ߴ
����1���^w���}1��v�4��!2��2��GY:_���`
�-Ǻ?X�� bK]�I��ǯ?5���Rp�TH��Ovf��L�ܕ�(i�-H�}�tq�k��3k�����?��3�1,S�.Sru���~8��F�|,s����NK*����9��qie����ܒe�垜�S��x��u{��fާ[4`�?KH��r�3J�7}�Ys/.3]��d�ɾ�'�~�������랐gJ�l����׬�:�S�ڴ�����K��61\��p5�A�Ok�(;�U�h%�����!'+4;f�8DHH���:mݖɿ����sy��d�ЇşL�0���A��s�v^�n1tΡ�z�k�{�9�N����jJW+�T�>Y�N����e�L�lj/��*u,
�vC+4�r�1��-�[;�,�z��<7��(#]����_.����F���c�.�Z�C�\$s'E
,�^�~S�(M$hm@9=��V>��1���|7v�븓� ���-r)�)�^Tڗ����T�ϟ��bǚt�96�m/+kXVI�-D�s.����}�<�B2[���p3�[�=x�W�~C�f�@c6-Ц��	jw�J�\��8B��
�O���FFp@�R�lFϰ�+��/f,�G��@Pc1-ba���|	Yz�kP��3�e��3��;���M{�,���?=O+�o��k2�)-��VB9*���GA�A\�B��� nPشm"?X�]�;fV��\��ҧ"&+��S㰞����{�l�?�]f��wPR���	i(�%8(�3y���m�$P^Zzp?#�b	�UY�����sӄ�����Ph���]������6u�\�����&��s��ӉE���M���M/���(>�u{�^����4�"H�ۜ�3������}D�o���+��,s[>^��4W�u ��#�ɲ*�Y"���b��Y~w9�l���6�>�|�	�#���̲���߭O�76{JBJ������+y�_�|��5��s�J͒��TN-!��)����_gcߙao�Q�X/�7��E�&�9���+iEfJ���MH��,�m�����Y"a����%g�'�fW.*"L^aG�&�p�B���5;�>P��` ��Qa���WT�b�8�H���m�v� �׫ z9G�W=��?������C9D8.��<�6_\�W�	���<'����!I~f���-��gVc���L
@�`��׼m�f���&����"�"l�ݦv�C*�o�{&�<&3D��;���.M��w;?�����:n[���%7 �ص�Q82�v��ċ��������j�˹nM��F��h�[\�!	��hc�=�r����@��BmI���+����Jk���r@���
����W]`�e����5��7X�\��`.�"��5Aϵ��j��J��F�t ����Ғuہ/�^{�F0W6�4����#�&�"��e�=���@0���y�%}x8E�K]������|����E��?>��n9���P[�=������>�7�vI&k��8��a�N=�b[�6�.Rh�@�p����i9��/�0���ϼ`z4ƞu���D����X\�ET6��=V���/M�P�n>uV��0���e�O�u�ad����������!��*[|Mf*,��u\l�n�s�	; ]��0�>�O�zE���4����va5J<C���I��-�4��a1D� Ů+��$�-5�Sg�W��Q�v��G�_w.��J��]�:�-�%�b��)�5]b��e;T=������N�z��O���{�,�����Q���`��>���
�^��rϰ������k�ar��U�sZ��I�;�u^r�+�;ɐ���cW�����t*���D�o9�U��e����{}�����4�: ���G���
Le�Y������D�x�Z⟑�1W�9��*��yTa��v(�����=L��Z�}���#D�D�S�ʢ�f��ʌ�L���*�96M��
��M_��8j����a_Rl�͛O����=Z[sF��Y�As_�۹:^�- ��7�O3��ء3�:�U3�Z�\%�_��vW���H/�ѧN���u*���B�
PC�q۟1����x�:"SqF.�s�qo�ܱ���i����j��a/�1ؤ��oqn��i_2а�}G�h�������.��3%�&1-���Y�	��)A�=��K�OK>����H{����S�?���r:�OŎ�_ ��ϲ?���f��@߀q̓���)��&�P��t5�<��U� qِY��ސ*��)!�/�fg�F��Q��3��j:�X�Ёv/0I$���Jjwl����ߡ2+�֙Rr��3a�ow�5JǇ�
c�>rF��9�	�Q�H�X�˶��^o�l{���r϶'���U�=�ei�p��S�7�b��x��_/��)g(�����pfh�� ĭy�ZvkV�
��3uc�dKB�@��!���V;*OD�-$t�-�P��仯�,3	�8Xş�b0�k�:J(�y�Va��;Z%Q��������J�B��|W-������RfK�^���t�K}a�6���w�]b�h�! �^}4E�'�ܗb��Lu���*����L�ӌ��<e|c���ȼ�g������w�Xlfx;֐>���_¡�k�klS�+��:y��L���V���n:�s֗=���U������#��W؛+iit����X"�����7�-�չ����^YםQ��'`�dȶ�y��2�b�/�!�e�Pb�ן�ސ2C꜇�^#uu�,��1�lS���F������f����wy��X�$e��������_Ei�M-�؍�,9�b�s�U��%О����V��J\�{f����1o��ˋ  ld ��2+�U��P?]���ac���$+h �q�������,��"ڋĞ�n�}1c��?,�z*|׵�1L:v���&���!��Q�cjG�?m`���!oȠ�)NF�՟d���V���_䁢��c��(�j�^������84��~�v���������^����.|})� L��(J��B�޴2B޳ ;�$���z�<S,��`����f*Y�Z!|u��f"�61�C��E�1����Y>��3 �+󑤘g�m��o�;��30Aӎ��X�3�]4/{[cV����c	���X���zK�_����>Y�g)ѫ��	P9[�Ϯ�I�!-�?럸-�������d<��B2�-A��<���ZЏ677ǂ���t�[�1o���l:���+厹�x�rA��3:LK9� K�ޯ{�/A��Wg��C���� C7�҈��iњw�)�/oG�.w~�#N�[��෈,_ߠȨ�a��I����V6�����4�&�E��y��������o���.a���]94���h�ӿ����۽G��r���6E>���oK���PK   ��WǆO2K 9X /   images/83b09b1d-e584-4d9e-8c7e-ad4061c788ce.png\{T�m-  ��)ݠ���(Jww��)1t��� ��twH7�Hw3p�������w�`X0�<�����{ވwo�1(0��j�t�6�P���4{�����*ƨv���Ro���0LQ���.
��/B�O�8����BE�����A��,����'^����E�=f�Ք�}��Jx$�&�����_��{����	����:�:��z��	�=�e.Xz���Ո^��HT���d��X�e4?qӜB��6���Ĳ܍uN��i<W̱s)���n+JJ��|�����H>���W��7.���,cr�����!������jS?m����߂�yW\ɇ���oq�+-���Aϗa�k�?�����wh����E���W<��R��\�� �-�}����o�o(s7j!��n�9��;��y�km~I��o*F�]��������
^_-9�\������t�{���H�Sg0JEQ�U�t�X*�oY{������w��ݶwO�j��9H�`�Gۑ~�����0\ڜ�۝\�J�vt�tƦ���Y���s�,���87�Ȟ���8ԯ�$���b����^���9��xas����	�A�)O&��H��s\OU�S0�i
��v�~��[�rԲ�����~��}�S���ʇ�f��澅���-?�+���o��]�S����!��7]Q�JWΊ����M̍���'����/�Aq�c���@�'b���bh%W�d��1¹�j����l�˵!mS���+���bZC�J�]�����v5����H�����/��J�f?	�gl�72.a���}S�ʢ��K�C�	_�=��g�aS����] ���ۘ���=��8�������>��x(��`ə�`�;� ���ظ2�$~|յ��[(Apy�
L�	-#�BM��&}c�6�t�����e-ݝ�>�r�mg����`���v��:ǧHt+�y�����B��[���{�ǐ#Eo'�(�d�>�YFg�Z��|��Zv�o6���v�E��\w����Q��!���l���u��p�iݨ��(���w����UԜ�E��791���V4~B��9a�~��sn�]Q?�͵�_L�{��{ָ{/S��^���25[�z��B��H��#֜�^�����i�8l�b�7���<��������d]�gl;�*ϻ~-�b�TN}�z��|��ӭ~m?�5�+J��jcӈ5�%��/O�r3oYM3�˰dL�z���Q�٦G�����v�8���nQ����'�`�η��u�4COW �O��F���%�d�Y^{\�#��@�3��Lݣ��8�*���g��d�p���vI�����l�席e�}\���#P�َ��+�6}��T�-A�C=�)�l�v��%@h��Z��<���aӚ�mwv3'ݥ*���|�������۳�����\����R}������	���h����P���a��_ss����̪9���i!U� qU�F�Q��]�x��|���tF^�4jya�)�jV�7IU����=�RV�`���)�Q#	~�W�K�?�?�1W$�,|a������r���re��-X$�Y��U��ͅ��<<�Hz���r8�Mʡ߈��T���������f�=I=\5�è�s�wP�|'aq�I�Y��/��kG��CH����÷ 
�lE�b"�e�E'��W�A�dF��ewŗ�@�V����~�Z���`|�T<N[+^-�j~�!	[� �E�'@��&���	5i�X�Ea�Z�:�����{���k��d4|�v޳<�oތ~Y��ƥvZ���G��Q���A���F??r��f�U���s�H��?����r�kA�2�K�|���ءs���q{ ����}b6(J�*�7#��a�˱���ȫ��TDC�D"�.��h��I83�Ŋ&�G L�ͥ6w��j;U���g�Z6�@�"����U�̩�p��6S��BjS
���@~2�t�����2Җ�1�R���T|������I�M�u��V��3�������n�0_,�J�j+꫟*C�[�
~\0.C��@���h��"ƪ8fdϩ��kƭާ��@9Z��Z�2��%���zUԎ�P*VE�s�gY���@Ŧ��W�'~ E!5q�sh��t���T�o�D��N��@oĤ��ԟv<���������}��DN�	�=owX(}�-`sAϲ#�zH���l�b�10��l��e��y�F����q�m�����`���� ���y��2 �q��c�Y�"�1���9⮛=�����I�~�3�U��-3﹮�(��Ҍ>{�a�A����ˁwՊ�(Ũ�׃,��5��F%ާ�ӿ9S�Z�D>#37ľE���Z7`�N�����Cz��D���%�a�Z�z���ruY���C�T���<B����!�7��ѣp�) 5�o�p���
ءEmim����O���(a8M]ə�;�E�������t�������a�@��M��#鼧 id���W�ъ���*�Q?�V+<�`�6.��i8ujr�2�����YZ;�}�lc̔��/���t�
� :��ϑu�P
i��)X�K! �����Tf�lϱ��Y(�L(��ȹ�p�W�Ⱦ(�����G��Y*.��#�-2x<�#��ǲ�<v�R�l�-ҝ�-�競1ԝ�Ls��gs���
��'��2�;X̓y6.�}���< YEI��b,�����`g�ݡ��ߝ��i��i?m�iww��Au�55>�R-�_/��D�e�k�将�^�I�u=��~c�,�N�EW��Ikg�[�=�����`\�2�����oY�5j)$5y��y��J�>���� l� ���q4�Z�(ؠ�oa6��q�1��!����kr�!|Ԩ�9�ںa	��*���4-_�̴������r�T��+�������K�Z%�)T&�x�T���f��e6��w�N�-������Fa�&�v
��������C�C���h�ޠ7�K�S���-(GА��`3煤���Z89�ڣ`%�	�۠�(����e��9
mr!#^���?�
8������"�N2*��z�48�okVٵ�� �R��;���K#5�_��tl���F%*K
>P[�$]c�ș������)���;��6����I�����v���8 :��� /��E�w���`�;A3����º��IV#��T�7�X��i�WVJv�e�[�x���|�|5)O�t�cfĒ���\i��3�uLd9��ދ{�W�1�؂�4���\��;-6��g̅>#�̥�a�[� uE����4�&��~�L�A����僨��Kw@l�U�4<ZE�5_�ڄ}W���y��$��?*϶vѺ�����p�F\z��N��'���rM�`�<2)����U��P%�Ի����-�WJ�<Fx��ܺnL��H\���ȓ���V�2S:�7�&��D%u��o3��@���Ń�~�F=�Q@9�&Lα�č慎ߙ�Ͻ^�M9����b)DRp6�R`5�~�@"��������Gk2o�9z�0�O�~�m^�����>��r,6[�3��C���#�c>���',�ʢ�5¬�h@�a%j����95��o�6x�d�l #���V��+v&7JP>~o��I�#�e���*G�2�������_o%�Q�~I,���V�JB&�]6�P�H88-7; �S�όcG��Q��������j
Ţ�mg�$��۱8��)�Ɏ D�����!�>T��~�����z9��rLk7W�-�x��BN�y�`�k1����7�
1er%F�7�h��F��UHbG��w��|��hw�T1�-ʒ�X�'�?p���r1%��]!�Ϙ���x�*���r7�d|����fPq�U�D�x����������tlW�����"����U%~�y�Se�4��)ؠ�%��%����B
�f��~A|�xA1PǎY�	��3i!g�r���xR�뽙(^MI���V_Li�Kw����E&�T}^����������ȼ�TW���n�Vhb������Z��
e9��vt�?Ò���^��q*���7+������Y#.h������8\�aEz��&	�T9���]����T���鑪L��4dz�1������-]*�s�f�����݊��I&�K8d�e<5>F�o�zj/**��G��"��jk�ƥ�V�^uDf��/?Kg�S�q	=,u0Ӓ��VV��Y��j<G����T���������Rjd�wU�[�y�p&� ���*b��U1�QO�:6�|~�L7!����F����5����D��dZVy�Cb�>5�ta� ��~�4x�� k�`~>}{����P������ǫ�S�e_N��Ms��Z���vO�ћ;a薓+�wzzy���Z�"���8tϾU�������KJ�@���wr�g5�Er���c_2�TsKc���<b;*!J��6��O�*�7��1t�{_��-$���~���x�%�K^�jk>�/�x�������yUz\Fvݎp�DK6���/Rc����X���{ޫO�%|!P��ѳ;&�2:�2���Pn�������N���;�P�°�Y47�m�Šʫ��2UEB{E��΋?DmJI�P(��S���	������)�=yZ�:��NĶЩ��Ɇ�_{���� 3y�;��V������j��H׀ܠ;.���(追�z��ݝ �5�q������}���ޞ��θ����_L@��	y�}w�C��(�d�1)�xK�y���'ꨶ�!u�&c �j���'�~<�|�r���w��2`��Pq�^Z����^��֒p�T��&2)�drw`�v��RUw��/���U�v�'6G��/�w`��b~�*sC�A�������)��d��d�
�~(�;*GLj�=�OR!ޗP�:xx�&P@ïq+s�D0!J�1���z�r�eȉ��<jQ l����p��NAd�m�j�L���ߠ�A�pG��x][>`�ί�_����[B���^�Ji�;��t�FA��[of�\����fo����L�ۭ��U�8�;����b���Ԝ��{D��ej�[��NXj�]].Q�q���љYˌ�h��ƫA�ͳ��!�<D:�r����:��3:��	GiVY���ٰo�^$=3�Yp��P9�����XF|X��>:��؍��TΖ�����i��R�2����1��P���L���^�@z]��FCz���祷M����%n�0�	���my_P/b���RD/r��ߜ���cc4qk�zZ�z���'��Ig�!t|��WA]�M cjʹ�
IH�˾�f���A������4tz ��-��a I��oxpk�1�Br�f����K�7��{����������3��V�pbKY(;4�Z��-�S�����O�Qd������+��e�1��v�8E���#*�v&Z���X߁�V?�]�6CE UFR�i��ɥ��r8YN�c�Xz����������a�Dy`�k2��8� �c�%%%4�=�E����ك��r~f�'�R+���J���*�L����('��0�dwi���\"�BUud0K�B�CB�Ѻ,
b��"�6I���s?�Յ��F�Wם�ɦq7PH/�սD5���lPXm��!K܂�%��	����	'�o��pJ�ʂ�D�e?�ل�,֍�G��(�\�ݔ��=L�����K�ԕ���X"�=�NFhp^��=�/��yV��Z_n�zq@?�[I鐅���@]�<x�Z�^73�i�.�(�X��;�[i�>i���K���
�m���I\����q�s�<Au'����]O�M[8^���,��� nn<q�7p��R[��d{��*F���J�;9��Wm�e'�J��Fư�h�:��˷�-2��ija6�e�Y�U�r����� ��@�:f4t�ᗑ��!�/a�6������uV���׆:�swZ��m=��A�@Y�jid��I[�}���w��t;����ho���J��$��i���
�}�F��6wK%�?'�����k~���z����c�)G��UL]Ub�&�""��@`�;� i�eP�|IO*w�����_ة4�g�n�����s����dLϾ|[���C�])
LX~`�7��q��_�>�C�=l�����6�"��`�$����%���VԀZԣB��_+���Te���l���'v@gRţ~���/�R�S�&� ՠ/D�GS�gJ:	�p/��H�F�o���P@���?\�TBz˛�|~o!N�2���>��I�������l�m �F�������'Z��)4�`�[08_�";�O*9�L6Y��;B@;)�G`�v���8���W39�,�2�5�UGL�j�~�zY���M�я}f]N1�'D{��}(k�&?��#�uuq��$#�)�i���<�]ə(�o�_L&����^VC�_�|W��a\���#9����J�g{D���%��7����`^tpab�ֈ�,��?�"<�<8�ƾO�Jk������0d�TK�Y�n˻�Y_	U`p�a�$5��le��nX^��:�>�S��Ol��ϝ�/{iUt��D:��=aZ����M�iY�鬝�;��g����2ѫ�r�AA�cY�pȘ�5��+�Zdc���@Т��4�͗<������zr���-�I�-���ｇ,����U@��&�|#��FՃ�	�c��֣3e�GQ��հ}���F+ANr����,T�Vm%K�:�L���eio�#v�lq���T�L>aK4��|#�O@�������� Jm�}�OO���v:g4t�I�U=�6?��O�l��)i%daP��:&WׁλTvƺ)��L���������b��!q�s������1*�P+F��X�O�(L���Zi���(/>J)ѱ=��v�Ā������:_�P4_E���B[(�nDN�3�StA�r�J��,oX��n�f���옫���Nt�&N��j�ˁ��x�M��C{���� t�N�r�j��g��ez����7_2=�h�h����\qܘ)o�q�`l`Ӵ�{����I2����+����wh����#�H� P>'b�A�d�3v+�A��U������b%f����L�R0[�whN��� s$�ϸ��x����cK]z �;n�Lm���v
��'ՋHӔ�V$)�P��揬�D�"�/��P9Z6Uvf�k�j��K��7���3��_ۨ��C$�7����=�YĒ�������yo=~Ʋ�Qv��?�)r��	� ��3I��^H��L��%�ν�B���fP��"����VB�JBz͙]!�<~��� }zR�Z?ɺx�z2�攫�⎃�w8h��@���W�E}e����l^�'�A��f{�]�`��6�Z�� �c��q�UR�o-^W���������6������t�G��{��16,މt�Q��O��a'e"q��V��Jy+�:��p;���w��P��;��YW�h(��?Kq��`7�
F{�6�#E@/O?*u��D�>�8xDQѲt*�T�������(I�Ĥp`F�:C�.D���F}z<������srJl��N��9�M0{��?d�����d<��Dݢ.�52���j�_w)�W�!9B�C�6�I�X'���5j�2�9#���&��[I�+��~[&���҉�(7e&K�c�U�uG��=��X\�pH<�5'�~�҇�5
v�`[6@h�(���n�s�|�4QV���K�J�����¹����"����\�v�	�h��X(��)��,�{	�LQL�!�l0��f��:���A@�i�3��xr,~	^�vd�-�:_�<�Dd��#K!1�{t����Rn�n����;���)������-��S�7�����S�X���}�۳<E�<��_I����5b���eMp�4x��'Zs��>����$d$��睤��!=��`�����8ʻ��t����y%L���@��k�Sf���f�u�wc�q]���ɓ]\'�l�B� �/b�w�Iڜ���A ���HW�d�E�k�/��%՞����әh�7`lj"'ߓ^婄�h(�S��yz$@���Cj ���	X�C�Q� �s7A&��8�Τ� M���w�6��]�MnyRR�t?�a����V�g���+���4����z2�H���#��g�J6&L��JX�ㄷ�V�Q_]:o<a�����h���C�Z��t������l(�$1���2��eR�R����D�^���\��ƐB�t�VIz�R���R�$H0��t[�z�Q��Bw���Yuf&��;����8�&|�#;�v��ޑ��x�3�Z���w�����Ex�%ѿsK��#�9�vZ�?�����:X�9I*⧯
)��?�G5d�˒��d5�_S�!�L�����]��r��)P%BOz��e�?��)�$�R����C!~Ͱ��<���Ƅ���Qs"�r/�7�G�&�/�)�x3�o{3v�7��wF�N�%�F�^�g.��br��� ���_�A�cC�����%�}�E[����W�Ç�k�G�����|J�^h�^�e	X��Ɇ}�A���������4���\��f���lD��/�����yK�1BكW��❾𮣨�Q�X!RF���oVT@�,�����c<�k�׸0���/�ZO�&���ۉ~�]ä�����eJ6/
4�� ظV.��K�N\4�������*��!���Dt���T׏
�-� ��)zP�i�2�p���`�j��֫�y����4�_����V�C�\����wj�t��{��3Z�ղ'��P�P��pa�|�����N�k���I]U|��~���*��m��g;�?Vg�3s�\��8Fx�oŏ=��fwk�U��f@��^�H��mŊ2��/-�|�1}����n���#�-8���M�٠h�e�[�����p_�0�h ��*Q"в}�d��:6c�[i%�NT�3�ɫ�%�E���R�I�����a|��³κ	��L� �u�x����)K�S���+:7<���>������_�}xC�B\�_��G�O-�y�Zփ1��!�(���3An���� G�r�h���ϫ{�_y����:di����7������s	u�صn���I��F�B|�,���ND3��e���)��͆r��Q�+Ƃ�;Y�I=&�+[by��Ï�bvjw��i��G��������?^��9j9�q?���,RN�2/+����-�;x��������Fߢ��k�p�YA�[P����}~�"f�V2��b2}<���PIs��'�)|Z��a5�)te�~R�Ql�N�(�B=�`��(�v��&�:�Hr� �g��߸����c��eRM�I�U�I�zӍ���ι��A>U�-���sF�}��dΏ_[<͹ZO�x���ҫ(̃�F��W���/�f�~����k��J��s1�y�^r�~W��!�\��Zܗ���e5�I���Fܸ���=ֈ?��Ui��&�$J��v��Wl�MT�RL�܊�<��ҵΖ��+�<�,����0�Ȝ>�W�2&1]�{}t8��(~�Cx��C��0<�Q�T�9� ����lreQ�du���$�c��q~��g�"���Z��Z�����,���pά���>+�������ք��\�|��W�0�2��$k=�$9��9���t�]W%,%�7�˲�@��3䠝�Nr����nƮ!4P;�}ANE��L-����1�Z(l��k�V#l���~}����^[0\� *�I'K���c�X�hc���Ҋ�V����! ��������2�����.��s�\����+X��[�<��؝�s���k�[??^*��}O��z���D��W�Pk��t���>�Tp[r�}���3�2�p���Ո&	�K����[ 1�sc��؄
k�tג��fO�3��E3">=�i?9�'~y�b
������y0o�����o<J^���L��N��X_G�o�0�@�<4��j/�P�dO,�c��� 7]�&�~�5��H�\
�c �C4e��:Y���}@��H�1E���5���tK�1qnA=���v
6)�0F e�-̰�p����E'R��`H.o���w�>2��X��8���s��8�V���_�=��w���I����N�U��w�N�[��ǟ׫�/ԋ�|�Jz�H[&�[vrV3�CH�g=Li��^3)�Zղ�7Y01w5��ؑf;`�� ��%�{9{J��˿L>���f3
�>��g$�\���zǀ���P,�ʳ;�������>�V��$�^�FH�|�O*�H2�?�z�cx�>j��3���^�jA	��:���c�A� �!M5�����+�m�R��(�s�������/#ZLP�ɂ��y��
5)*�e�q�	��{�(2����R�5C�4�&�H���)Bxe���1|�O�� /!��[Ii��Pl�O?ɤ�K���0_;;��jA���؛�Kފ����^.�#&��ȴ�#��,�f��Lk`��1)�~	?%�z�� ����O1�['F��i���� �Z���Q���Hv�����XUE6;����S���HN-��}�BU����8��E+�����c���������n�\�Db�
���$�{����ʈ�Ѓ'�ج�o��U)E�I�0�2Im3��c a�h.T9��s6A�]7㲁����h3�Ao�����r=�>qu����[���/H]G��\�{�ٸ\�X\�P�OJ1�*JA;�C���82��!؝�=�G­JQ�V��PLR�ᱤAS��`�5�>�n�Ŏb�������޼�:j�ƕ�tŹv��	���Z����qj����H[�`kEv�����t$T�ٵîJE���]��~��N���i�����Q���|����1��n;v��Η/�#i�������q���S�;����;ꋕ/�
�_�5I�x����ܨ�.�P-\�̹
Y6ݎi+:4�T7��]f�U�T��N�7fC�!)������Hi�|A��,�6�_�+8ܚa�N���@��,^G���s��y���Z�u1�AZgc�V��eW ��g��t���Bl��F���o϶ǹ��j������M趒�f6�����/��۟����.�Z�~<�y���h�wJ��P`F�|s�kM��ϲׁF���elM�K:c���A������/c� ����>��c�Jr�K�s�rN(�W�zw�0�H%cj5z;�?�P��OP����.��X��aCi{f�H��%r��ճ� ��hhU�$�
�!�慁�g�J
:���T'&�|�#[�2�'%cV:ŧO��/�i���3��`X����J�+���6�J�����"T����-̸}\��Wm�|���g��zJ�{�4�������l�k��QRrc������T*O�3�UEEE[�� 
�����^��5�Јd\�R_�i%�c61D��QE&B���!�O���x�3!�W����I���qɿ��[� ��7��7Z����U��r�iڃ����;�ҩ2���г��㊆ZF�^�G�{�	A���<){"�D�����O.vx3�m��F��Ɠ�v�Q�z*�:��M��v��:fi]qd0��^֣��v;�y����.y�,4�O�@o{���Y�ʏɢ:�}w|(�d&q�KG�:�:������̘y-���c a�<n��%N�+���i��(+{`�5m���;|l�^�������u(��ncF�T�4j	�.���,��D'�Uh����[�ײk�/ ew2�(L��2?��^-�HH�ۉ,c5w�bʿ�����3oQ�� %�q�<!9|�	*��u9��l�k%�Kk>��xy���iH�IM�/�����*�D���OϽ�+�H�l����������9-���֣��%9�����v����;��4	�T�����Qx�X���'��?�[Ƥ��jjPWjJx�v��3��˸��|֓Jr�$�w�kť�(Y���P�y�nK0�3 �ٍpڣ���=��K �#1��G��տ�X]?��?T.Y?V���X
s��t{<�:5 Ī�[a��|�y=����[�xmJ��|�א�`�f䫰�롲�!EE�Pp
w�Y(�2~�@ ��@K��VZ-f���0�ލ �Rǘ%�)bQ���,�a���K�<9�E�y���h_���|AO�,�M��z�.�<M?~�P6��Y�_��B��{�n������0�ƃ�	D��c�� �F��ה6�^�D.8��cPy��"[�����#p%A�Od�Ƀw� K�y�BAS��{�s����9���;��p%��"����M�LҺ�z�Y���&�\���ZC:)Q�H�mU �f�@���8�qp�2���(tc���((tH�n�~�����ފ�5^�q ��M��!�W�p<]�X,�P j0�%p��i�X��4���+��f;�YU�]�K+-)!iTf���+�?7�
-q�,dtr�x�~A���� ��'������qk���އ<�a^<�u?,��q�ߦ׏���W��^�)�o�k��A��PU�=��mߩ�H����۲���-�)���0�,Q��)�{��<�w��Z�%�Ma� L�B'�n��di�<�e��y�<�e�^�Yno؃�u?l*���o��VWl��~���1��zP�Ys������p�x��s�%��S�:����֐�W	�m�^#{���b�MG
t�K�\���q9�f=_xp�lT	i��voF�@E2q�*8�� ��0������p�&_��1A�D����eK�J���ӟ_�Յ�yL��	Y�B�e��a}�ݯI���.�Q���M6���O��P:�f�d��u�Pd5e�جJ@ %��7N
.���}5�m2[�:����uC��ώ��U��gL|�oH��I�����?&!M�]��`�j�L2(e�>�v{�yxX%��S��m�������g��?�w��~nŊ���5J��֕�r�ͪ���K�n���]ש�����{=%�>^����D�&��p�V7^���矁 ���΀�ŜV1�=\5�����9��˺�{���$��b�*���d��j�h�	4ڊ1R�L�������^��#�-�jFs��V�e�|���#�;DY�o�9pr�p��'��&�{�%�|4���V����W��������j�q(���u�J����wj�v�#"l�ڙ�7@&a�
R�<�����}#���p��'hn6k��CEj�z�\���;�|���)/���H)z�[�GE���T�Q�]���겲9y��V[�
�#��:M�&��C0O�>�*w#ֻq�b-�đ��]ok�?�P�gϔu�b�`��'F�?�N�w�AϞ��>�:)�A��V���CC��~�aǇ�aJ����@i;w��d����~R��Ճ��#��({3�h'FxU�`V�Y������S�����~��ek%2x(!�͓!�ypBP��0=�
�;�m #�ZW^���^�3�j*�G�*c,f,/O�p�@���(Φ���m39���Q�G��j�t��;�zC��Љ#y�5���r���Ʋn�N����*~��6.~m0�F��/o{^1AЇ��X�c�.=�:���vZ �)�pK������Xy3��켴���ׯ_M��ތlY�8�X�2���.{�82o09r�:���!KBLcc|��&�#@?���E�)�j��PZִ2��j�<� C��9�_�(/~v ��
5�g
���h���=���R)%�U�{��h�65c��l��Q���U@}H4	�|B�VZE�����S��T欢�"��)����	���ॖ�v|r\|%�z���#�/�	�_�h~{8��ה����R�Bk��H���[���H5��RbD��גB{p�$�*���k	4�N떇���ݦ���������H4�(�C�
#4�~Ȓ\�FV�]�̭@�G/[�?&2Et �ӷ�f��jA�+=����Ͼ������N�+^�#U�^U���/PHP����+Z�^]warsd	�φ[�4�74��5w��+����ePY��u�����Q��'�Ɂ�wˈ�h�����T���W!���i�+�$�I�{Al YMlt��o=��ڎ�C��ё�4��9��o���=��c��/|����~�ЋL(��bԕV5�:�S`���|�����{e��o�w�K�e�z�D��^?� ,�O�=�Z����R��|.%�G���VFܗպ��p�)�˨�K!�gIHd������R�y���֚����C�� ��ן�B�+�?z����t/���	B�`��GA�� �A�@�q��~��E���]FAX���5l7�����3���������������Rf���K'�v6��4��:�i͈�#��d[�W%�Z�c�':���G����FG�EӰf�"�3�盶>�3<u��>C��僡?��p �~�Z;,�����L�	?�蕱�ezD��X����U�P@zB������Snr����J���㷴����o0�!���U10�)���Қ@�C�Q�e��S��*��ȮoLtc�We��7�Ņ��9\��_��Xi�����������ï�=D��^�q[�v���ѷ���.38ʉ�1���Y�J�V�n���7=jXrrOFU�r��l��W���ܭQ{����uK�O��Μ�s�v�N�_%l�!E�����|�_V[�KƳ�Ijd�o&,S����=�����H�	�\�I���z��Z����wH���_��k�I�k�/
Lҝed�֝t
����I���-�^�hmG���IKGް��+O�؏�d��l ��"�~7ɯnF�����ͣ2oA��$4�{��[�Ib	i�$� s��Ϸä�7��U���bR���7If����++���f��df�8�;��S�"��eR̬\B97;i��>����n26�U%au���q"��B(��gIR�B<��pj��
�p��O����hζN��WU:�'�ꛙp�� �zK#���!��P��-�k�v�ۣ��ƛ@_G~��=�������6�[@��m����G�i!�k��Ү����/"���Q�P�pmy&CiQ�Ƀ#�d��~����L!���`��+L�A�ji�8�ݓ� -����唥���מB��4-?��a�8��s�#v��3�&��ŋ��E�%[���i0�#��T1�i�z��5&ɗsc�mw��=o�(ռ~� =�oX�5�\��C/�1���a�����s}�+���1?j_<ޚ��u���^���64�D� ��ń�s)��80�)ג �\��7F�����H)V(ӈά�����4��H5���y�φQ���e��]��;+�;�bX�E)|H��')jڊ6�d���9�C�Vp����:�%L��8��H����Ԗ�O�ev�����g61!Z/�l �bOŸ�n�Kgʓ]�Rn#�@Bi���%P$c^��%�q���:.���բ�XH
�^MZ]��}�(D°�k:1�[]������=�r#?�09�
*�;�G#0�j��T?ت����Q�d���m�G6���5�q��i���u��T	���g�`'�!�צ�.��
񼌔$��Pb�.�������"x/Ue̔@JHC�o�k�?3f!�c� G+|���Ɨ��nߦ�@���.AD��چwޛޓNC�~Ս"�GS}
�D��Hț)K�K���3*}�j���vh�8/`�J@�ދ4'���p�?����R_q��.	�8�XtBf�ϒ����yn�t��Ɉ�j�rn�vu��d���V@�4�n-�o.�eXXx��CšTF+KJ�Կr���\�3�%�b��P����FG�F��f��"�"��*c�U�3��>殐,G�����	Nf����T4��M��G��Fem�4٤�爊a�=���ഞ��bsg�#���P�#�#��d�vTy���3��%�Z%�:�޾���%5-&��Sg���p�X�`#'��G�xz�7*��2q�r����o���=��h��>킷��М���>Xv-������{�͞ܥ�Z�{��ko�{HgU����X�}t�R��7�O�}���ߌ��k�D��3#0�D��SA�]I��]-YIG� m`rץ�9�"���ߚ�8X#X-�=`i�d,Q�M���Ua�S7���j��1�Ǝu��&-�P���Ʋ�D�����!E�b���{$�1��=D�Ыn�ju���',*��
絶#��������u*��Դ��i����d��amj��y�/�r�X�^ߎ�wri��o*X�:��=�e�qΝZO�|�c��K�ED��-�䟅��"�S�H�w#�Q��+qCg�@({�7I%R4�r�ア�#N���u$7U�h!K�׳�T!hŧ�UMa�A/�,ozt����1ܦ���L"���%p����G�cG����b�l��\��-��Yx9R�Mt��~j ���VV�@�����Z!V���������{C�o��ه|=	8z���:U�?����	�Ln��h��f%Z�=�+�c��|����T��� :H�=�p#�u>*<�7Y��tձV��[@���O9����s�?nn��T����`����t�x
(b���`:!M���q�[�riD1\(��>��yH��A!�[�p�p,����#��%�Et{�q�1��ܿ�O_�d۾M���6��VAb��A�Q*��`0�K$DJ-Hw��*-"!%����}��_�y]��y\��|�	.ѳ�����3�7�d�v7$�ФIF3<�o��]n��&��9�W�?��䧪�+�0l���u:���YǟI/�g]`KN��J��p����c_��9���[;��]*~���8���r�H��j��X�
���3x�`0�������gw�\��I��f=�n��r/����9��EL�,v�@sF���a�vz�M�dl��#V�����Ѣ�s%��+�V�?J��e���~�@SHKB�R����8�D��P��������#В����Z9˙ݳ�-D���,��L�n*��������Zmh=:�f�V7�t}������/���-�E���mȫ��<�~-��.�1���v��q�{���Y
~�Nr3}�]�_��拽�����%�3���B�o������c�������DiD�=��Fc���,�d�Wc�zhGC����_��]�KS��.8T�ʏp^�F<����������0n=�GN3U�^��=����F�[�M�`5��l�;M��|4*?3��9�mk"@I�
�`�p�iY���nW�GL��m��ޗں�r�Ĥ���[y��b!��_�L�ٷ��4+��ow��N���a��j<����4Y�;Yo��c�����%���&���}�A��s,w�'��gHb�p}����>� Ѧ� =$�s���eԦD�,�QO���_��"��̒�(v?T�Z�L�JQ��4i��Ïb���m��d�yO@�F<�[�C����	]�_�T���P]hJU��R75/���4���$���늬�ڡW�~�u��9Ϝ��K�vh3C�Z����c��aWw���Iؼ������ME��yϹ/Ui�C��?Mk�y����}ϒr���v���=�Ւ���5��Ɔ�����5xwu~���)/�o4ǻ��f��$Q��В���d�x�(|ZT�a�cU���z��(j�G�E�,�k���))j�p�6 �%<�r��L���k�m]5j���h
{�)��0,�5O��y�h�U�S�;I��K���c�?m����:�����2��!����Q������.��=�b��𹏀|b��x3�+=��)�M��!@	ZPos��*H�g��շ�]��RG�ѷ���ʥ�D{�K�:F5xmX���!����L+�) �N�3�b3�Z΁q�c_���ӈ����k�	�ĊD�Έ}8Dw���8�O�ԑ�{�Y�;��W�I[�-S�G��F��0��\�|�"Ie8䬃Dc-�R�$N�v><vU���ۑD�����l��:��8�9���XU�G��a�8��?����(���
j�OEz�m7�[�@���2Six������|RV#�ve@�y򲛾���{s4�A�\6g�ߴ��G~��D���PR�N���r�^�����r
��W����X�:U�Y������1�������?m$C&����.���;C�h]��T�"�=(�<������?��^SAp��<}"�Z4��0Ц&n���W�ӶEn��A����Q>?_�:�]tHOU���$2s�,5>�"�]
�$w�ڮS��߿Z7��rx�c����;���0nBK������x@{��AL����Ί�LV�9�c���]o}*\%���o&��*,k��#���@J�6 %u .E�n��4n)���t�tŀ7b�����i���ċo�I�
Pv"��7�Y�&���)z���e��&���6Z�������g]%V���9)הW���T�7L	�һٺ�*�~�4���wW�E�U��%*lż�ʟL!(�Q_:_����{]8�h�G�C3������T��%_%��������'��$�у�N��+�|���n�Nwf�sAw*w%����qf3���M$I�:�))��������]�>�$�)�N��QU�m��� IZ+}�\v���~Z�=�鮘l+��pF�W! ����R�T���t�>v�z� 9I��X�'���/8�E>�2?�U��=р�]�5�w6:���)���q���������:��_��/�(��Q��������p��P��k؃8Ħ^s�!}Tw�~g�qC��&l��/g�ӫI���8�
���j����5��o�9���p�/��A@�~���:ڿs2�8+�u�0��$5Q��ׇ�#[�[,ܤ}6���v��{�0C�����rB�JH�˥�OAH��\�7�5��X�ZE�PG��=�?��>1*9��m����!M�,�	3t��F6�s�E�������ۇ���nyT$Еu�<���a�gd.آN�,�5���q�%*��@{+��m�Yoz�5��ο�����
�
?������������6N�,�4��Wev�M�W[�"^�^Ld9���t:�ݦg'Mr������B.
<��
�����K�x?���̼��Z]ߙXW�Ad�C��*����}=��N^w	�+��!@'����f?۪(��"\B�V������;��V���8���d�@~��j�]�� �%��} �l���s5�,��wf�(+��k6n6r��)�u]ߚ�u�hBA�ةP "�����-��
~{�	����m)�ݻ�,��v���`��
�9`d#�,�|���7��f�ph���<쭬��Go�x�P����@CB����=L>�*�!�B��a����'�z�v\���:"��,�g�a<Y�F�t����?>�c�ͧ?����ڶ����l�1翙�\�w���ct �������UC�k+�A��3�Y4�5�G�7�L\E�P��L��"�����n$r쨯��$�\�Tޡ�Lq�cާ�Fq�aH��..Y����e��)���Ͽ����Ӑٲ��,�o��F�qn=�]l4<�T�Mk�X}@K<������~�:���4��~:�o�B����Z��@�W/�N61�$L��Ĉ��Do�/&��e1�9�(	��F�>ńX�A�֬�z��L�'�ۓ1E����� ��9��f�<��T;&�ХԂ����t����ZwhV��� �-y�U)��`��?�<a��`nQ�'4���qoB��e����X?.n�����ea��?��V�Smv�}����R����ڥM�6�`y�|c;}5�FQ��	t� ��$�wc�W��ƃs3q�ײ|��l�_�,<vxܠ�D4oѼ�vʏ������� �8]����gHl��X���p�)R�1Q?�.�7�%
��o(��������b�)3Ƕ;��[�uuν�"����?'������S�B��
I��e���x�i������@枾���)�d�a�F�Li%����":�~"��&�9�[�/(9{�I�g��>ݺ-^q�b�V}Xk�f����tɲ��9�N��Bư���Ǽ� Q�&���s>���"�_.T"�v�@uHt��D6���3
S�#���(� s_<D�*�Äd�[7���-�݄O�|5���b�*|b||�����OЯ��J��vkgL�*N���U��J��V�����Nq�P�.�r���ÕV*i^C&
�X��ҧ�`�9��W��?E��>����E�?֢��m"�#�6���
���K��8œ��R��A'�~���x���NB��v�����U����RjcG���H"B��tg^��"�����Y �$u9����|~���Ԁ ���X��������,^��VMu�p�-�S�&ߡ��v�VƱ~�����zx�~3|;���W��0�e[����#��q*
yDśͮ�!�ӭ�R�v|+�Q��B=��� �zL�H�Ռ����B��-x�0)��O�wa{�Nu�E�I��	Ͷ_|���ْ�'�����%���LA0�ȯ��D;5ڧo���vMN�Ni�3&R�\vt<t\�}ϊ��,q�#3l�����t,2)��r���v�<j��*hH��r���qTUK�c�HT�~�������z��Z�#q���/�Đ���9� W�|� 5�??�C�h����߾��ayD�v��o�w9oJ��4	��${G+ޚ��v�,/�E�Iڣ���e��X��$>�z3|c8���]w���{���7�m�#���~���
$�K���F�������5���T76c&.i����b��Ƃ�S4���ƒ�v��F$ƖɨOn�0�h�� �"^���6��t:���V�f�'+m����f0�ˀ����V�?ʀ�y��y,+�lW_3[7W?���~���OB��_8%r�[M'2�J��Z<پ�t
�`a����a`G�-ޠ����Ax���|�I��w��I����{xd6�N6&�$�A4M,ES�g�A�@IM)պ��Έ hEX�������Af�wY�~邗��,�B�PJ�q��ɐ$�s6Ů�,Hɇp��;I�p#�_�U�'Wb,��٥��L[;i�X=(��n��ʜwG-�ȟ��s܎`w h�$�ِl@J��y��[3���t{�N���������J9��g�s��Fj�B߻��u]�8*g�X�uCKT�9_Q7�І������i��C�ҡ	g&��{�D����w9~_��� ڜP�QB�-94��E4����W��݉U��ӕ�;Η�Z�`�P����ՌF޿ Z�l� �hQ 1���#�jh�rlV9M@��������oQ�����	��~t�o_�.�LF���S�Ii 6�(E��YM{�)��<���-��V����0���2�#D;n�b(Pj0f�/�(ЂY~�)��~���±r�q���, 7���.ܝ%k���F�O�(^��:b��^zd��[�'�Kp�5L����j(�\�4�z3GƬ3dg��>k��J(�0f�88�Ţn�DD�3���O'�2Ύł���SL��pb�����8S%�[� ^�a4�'�ﵶ�����S奯*IK��;�9��ǋ>�.]��[�C�I�>���P�:�E�Z5�I��Ḥ7L�!%S�"Nf�Cupѝ���]���x��U�}���\ُ5�W��%���9��$�n�HE���d����Y��Q���%�~0���C�$�����^��'���o�����kȢŖ���|N���I��`���c�]���Tb�|Tn0R��,�`�#�[�Ϸ����IHX��񻟵��S�7��-���,��� ��o)�+���zL�@�B��|Е{�%1�W@�8�,�]�c����#R�y<�>zU��ӥ��:hy`:����H�0��5�s�UU�<�fgaL���S��7o?K�|��宫�d]��7�1��	M�҂�V���!��G��5��>���q۟���{��fl&���m]^z��zH�.y�}/��=.��7h/6K�Vf+�s�&R�j�� na�uZa���:~/6z�4!CN��3pi�.�x��x[����x�&�! �G�Fs�߱cO�T�>�#�Da+\Œ�jR���w�
�Iǚ�Q��K�x�Q��Հ��v���F	~��%��Om�^Yj�jͥ�2��/R�.rH�4�T��D��I���'��p=��j�1}��p1-���PR;x����DW�
�����x��/���$u�TnKFn�2��g�b�x}����p����g8��<�op�hv͛���y����V
��4�g[S���/��� 8���`��?[���;8��^AW��V���W�G���?��r��^+�o�jp�'B?\��PͮD%ȧ�L�j<����)i�T�"t�P~�Lf|&@3�㥋z�nQ{��,Sڧ�`hiӫs�C�[�D5��fu�)#EO�QZ�[jċĀ5Tl���B����f]���Us�Jћp*͙ݕ|�4����'�k�ju���R��Dx����t�)��t��;n��XR���c�׶<�n\�V�M���� �l��;}�V�[ٍ?p#�����`��_�dV[�w����7�}�;C?�?S�����}�����D��y.�}%L�&��S�]���qݯe}'l5X��u������xoJO��92*�iHB��#s(U[i�(
�����r�(�tكy�h��v fD��i5bN��C>���uB���Ră��Ù�c�������!��O��8RVAC�U�=~�é��(LD""�%��$]��럶*t7�/o�8�J￥���:"��=����	�����R�����g+
��V��W>�R�r�KrUi�)OK_T�n�F�e�8��,���2�8X ֯�C"��W�NM?�z����p~|��w���x�˖?Y�����w��$�%�_Jo��մ���-���9u����'�
��(���w�5�1��6Zt@.,�������vkB��G�J��
��t�,��	)ܳ.hY�	�<d=1 ��ɯS��8ra�Vxޕ�HTJ�$L?�]��*xC)�m��Ij�&�v t��D�l�,�Sx?�l�ݓ��Z��>uR�b��h���o��e �E�>����i�Q���5N�՞*���dMU��/�&V���5���E8�c+Z#@����(}ЩZ�{���c��ZvGff�SIK�����h�@�u`���ͫ�w�ǲ�>����9T���~���-j�����.o�/������*�;���~q.t���L�Aw$��tD��2и٨6!�|#V�����|uH�jD�F�B�}#�|F�"��$�h�L�OU��I5�gx\��T��A����b��"z�V"V$ۡ����-���vV��ǋ�^�l�$�����J�"ɽ��l�|p&R'�:�v<<}'.�Օ�8h��EpU���f0�i�}���dN�hdm����$�W{��d����h���/�o��KuY�g��
���>�S��8������A��X���]/�j1~N��Rx� Z��z��ź��E�b��.�/�<��5�yAFRr�۶X��h{�Y-ˎ������ ϫ�\^��G�2١�c���v+��D��ǎ}�^��{x5��"������5/_�����U�s���cC����03AR��z���c����&����nKOg��)@}�����Uaz�Ȝ�	�'$,&o��X���$\,�a(��^�^ٳ]���p�d���E}g� �GܧS��c׾��tF�˧�~h�����1Jb8��3tM�UEmAE�ˡ
	�T:�Nj�M=�a8�r�q�M���#�'rM����o���^H�f�s�U}���>��)d��7Z��v'�=P�`W0H�{v���U���y^C�rWÁ��=�Ț���,1g�ؚ���o-+�3U��aiU��%��Ǒ:H�>�#����X���L����}6��n��ӧy2{������d���/�W��Y�~F];��ʑ���˶.^��x��v/ ^�k�Y<c8[����߅��3Δ���u��~kxO��"OID��PV LQ���k����f���{Mk"X�oY�I^��*h��`�bC�W _��f
JXgn@���"6�
��Fr9�Fv��Q�RG��o�|w�� �ۼk�0�*�.y���h�"���h*X�4���E�=�Z�f^m��XL��w��F�e�H-� A�#�k���)���#2�q�m�Sg ��X�vC��,��N�yZ�
S�۸�����_�8�>�5�����c�<2&u/�t�f��	6�B��P`�F&m��[G��u٦�)�W?�D�h��mot��w������t/x<W7t��v>���_61��ONNKO��|8C<Ǚaap_�?݋9�����+������_^ng ���PdNҵa���a�)*�t���fe���q�)�Ô�U�h�èf�>4��fI�g���n����1w"r�)"8�t���]���=�B�ԏ������������5���D��_Ff�#��(���줳�
t�A��SQ+�9!��I�����	{sw�Q���]/��^�K��T��S���m�Y��v���$Rߟ�
,�`3Z�$i��j>��]������'[zy�~�a8amǬ���&'����A�Ŵ2�jC�>*q�T�g��$� j-��R;%��H(U#N�棆YM�'s[�S������_LUe%g^�r�(�y8nث܌����\��C��~�<���˔����������ڡ�.��jc;��j�����F�e�?2��>�����q���&%N�3Xv��P	ܹp���}���%�[_���QWM�T��;��a�a�����^Y��~���/A�"����K��w�U��_@cFw��4�0��8}����U�fOu;�`8#��~`���nM�j"�y~}zu����b'�:�Ĩ���rnSM�NU=�u�c���c ����;bЦK}s���6���I�G��0w�R��o������8�>Z�(��!k�A�eAh��Z�����H���߲x(Ĳ����f�|���à���]�"1� �%�J�pKT�l�Ldf����U����\�}E�軹�.�j���g���󮬬���9�w��Zv�6�<e��I�w�7ǿ�ܷ��f��B-�	����J�����gn=������Z�:�'��f�x��j�f_\a��u���%�{R��M�ӀM�����4�6b�QC�u�z5�e��rd�[{~:J��#ɵ�����y�#�%Y�ư�%�<;�	��R��S
�(�X��rj����N��~---��_�7;ZB�m�ۣ�,�gB�=��1��87G��{��Mɋ����Tx�\�+WC�v��:)q̡L�:��%P���1��!�ݩ���/�Zh�����������!��;�p���t���OOq��R~y	S-��e\(�?���͐R�lu��<�����ƭ%2O�,~>Ҩ��n�~a���i���e�Up�o�0-��v�/�6Wޟ9����!�������G�dhUZ�nl�Ý�dtUa���A(�N�?#�$�U��IME���I��W4Tgtb�DHJ,�E�Z`E�o�1���� i�h��t�-}v�,��1�i�}��A�T�E�C���I�N��,|j𘓩�an��&��E�)�.	u"m9V(��\�1�����(�ij^"��BD�d���-(���ٗ�ՠ�>��`�����~ ����H���c/�	���s8�����и��w׳o��ց
a�x@�����l�3�7�A���@〖㩹�:�l#S��F	�3_ؽTx����qmT�����}ר֭'�!������=y��ػ�,���ףc���R����I-ɀ����;�'j��sY�p�r��=�#!	�qa!3�PdHd��a��;#oy�-
/VE��8��jg�����aI��G[�[Ҫ{T��4;�j>��}��jtZ>]�gJebq9D(d<ɮ�ux�H����KI�j��2��P�,ʥ�r6�#���@��*.�&���k2��<#�p�z��;��6��]<O�-�c��x0��n����~�L������O�iU"�v ��c9O}�)e�i��$�9&��Ѝs�~§Gh�nI%^�8]$A��\O9;�4���S�tӲ�3́k�^���0*M8�Ѳ3'����Н��/��3%ד��*�ʞ��<��&�_������pë�|'�g��9��V��筧<���m����Bz6+=>eI�IG�@
_Ai*)��",���ÌVc��E��)�����ZYT>u�H�ς�m�*�������<5X��ȸ�8��X:1�SCUR�9$�-�<��#v*m�rb��=B����WO�'������f�Ǒ�98j�G�"Ζ9�� �o�5��#&U��L�Pr��=���&#�~xY��\�yh�u�|�N������*�wg�jLz�ΰ� ;���fpE�-u�T߮1v=�X���Л뻷����6��ʬ�*�"!�ɽ�L���w�1�w?`.�W%��)q%��B���Yļ�gG���E��!�<���G(�������}�w7Ҝ�.Nr��a:Y�启i�ֽ��4�W��߿�k�G�����,�~Tna�6g�udֲ�O�Ig� v[�F���M���mEbk�D�Q�6+j:D����k��m�5���P��|H��S������R����-�x-k�ҭ�.]g3տ)}������!�����<"ꂪՋ�E���`(Iؔ���pXk}-�%"��:`�@�v��;��a��j�p��I���A��Щ�k�i<���	8��lSAV6
_��8*�D]��e�^Z�鹦��質n������cw����O=���W �U|������>�Sy��D��jy\̊v7s_�J���6���E�iH�WC�����H���R�J��S������#�k���H�����w0��j��5=SK,���c�Bw��������ث0jG���	O�Ƹ�T����[ʘ�"���U���(B�5��D����{��?{_G��ع��K\%��V�Ķ�}3t/M+�ͼ�1���,���S�8Us�c�c����*�
�R�Wb%��dyC�?�����pi�r�(������|!@�ȨA��]��8���3�yﳾ��6�V��1�/� ��W$}5�FʙHϽE�f�m/9�h|�a�M�[��~���07���o`0�����ø?����A6w2N�z{h/å�[��\����>���}}05?O�s!��4=JN;�l�p�1?Q^Ꜫ���K~�0�'Z��ss���Ik>�eE$�լ(�U��ܒZ��F��t0�R���c��&��{+K<��z
/(ȥ��JT�9j�PL������p)K��%�F
�R��������T6\J���[�c9��i��_D�ψ����C&�(�y<����l(%�Y�}L��QJ�y�j{�I��`��X��MvG}�$�^?���J ����(HazT�ѷNA�@���mi��L:������ٓ��>�ـ|m�X|����퓿�C�����Wԟ�w���hH?b�q�<nu{�F4�1ߣRkٲ�v��=a,��|�]`W˲}�E@L�`k���.Y�$�{/~�
ԝ�-��q(M�}vf&�)H�����^M?�޻{� -O�h!G\�ܸ���nly+���e �6����c ����N�5�Zax�20n1�x��vW�K�)� o0��F-��.��Oڬ7�z:�UZ�B�;t��-X�Jr��P�\��$K�A?��?��쓥�g,����O����x\�h�CE���C��g���YO�H݁;O=hB=�,=�b�_V;��tK�ձ�NmG�7�W�I�F��j�$~��1M$���������A/[���E�`Y��U,H������iu�<��Y�I��<�gU�GV�~^!"����&��e�U�x&��$������U��u��J!���څ����1�&\�'Փ�?��;+���=x�>S�/(���P=��_�Vu#X��:Ӛ�������P������!}���[��,]�\*�����{�٧����{��"QXl���S&�Rm���q�����kd{[Dx��L�D�K#K1;+���#�r��\��q��F�.�cݛjK��t���E���� GN��S]�GlMܝ���x��{H�V����H����Nq����oX�C�d�H����J��e�誺��J�O���_l�����+-3��n�������{�!���#�:I	��w3���.�*���0 ��Z�ħ�56���^����p�Y�x�����DB���_Ȇ�����\0����厰��.��'1)?�\�I��|�˗W#�y�mWc��C�Y�m���E�* a0TXA� \���h28��i5�O͆ه"� ~Ko a�e���Nk
���)���N\�����R#��y#����ǘX�Y6���@h|9�������6\�.�pS*f���. r9*=�(Ԃ�w(�KgrX��W�8H�N�y��/c�! ��N�e�����dW�T��qV�-c)԰)����-{�i�5����������c�^�0�0ůg78�Jedck��ߴ<���h%�O���G���/�����Rț�����'ȻGY���Ō�,�d��#��Fu~G������ݑ�M��m�n�H:Ϥ���Z巊>��S�	�*R`y������i�E�QLt�\�0X@�B�ۚP]4���~#�����h�U`���6u�=7�����)!��S���2���+�"_�K�z#��ny���<�aQLv�����������%�zuW�w���f��auY���v7m�R�Sk"E/�� ��X���)�*jDl5��@49ΗrZg���\�//���}������Lwl�T��jIN7��B�XC������Bzo��U?�c��Ο*�up���W{c�%�*�}�ԃ{�[n�T��I2��<���e�
9
�B� ��d��v+b޷h�����1hUћ*`���bkJ�2,A>p�s�<Ǣ�eӴ�5QSUU�H5fljj:��KHU�Ɩ��p��jr:4x�
`U�} ��`
^�9 ��˺�x�JO�'ik�[���Ek�m�*OȘ�	_i�5���`'+G�C6���E�l^|	�h���?��P���n�Z,u,�/]��H0��L��Z��oV)u|1�!,i�Ks��<�����h+�k�uе���TH>�����Q�`n�1�`�qTV1\�����������]�5���"�$s��1|��lH��(��_%��m_���3[6rd*�T��=��z���%��{F䃣��\�W�Q��?}ײ�E�z����b҈:�,{;ՠ����d���v�;.�w���Q�i����]��/��'��}���VR��~���!�0�* {��������zD-J�&�͂Jj�k2՝��N&�M�^D�<'�>Z=�v?�%��AE�+H����W�޽,f���$����Ǭ����&�3$a��N9I@[��:��z>i��~o:ρ�}��E�{��^��T�P*�ܝ��f���6
���d�:q+q\}�����H���$u��}V�s�1~�'N� f}܇���t@�^��t�����C)�/t��>[���1?rz���c��=�����!���_�G��D�)�_�n��j��Lg�Cq��,M1�<���eM
�f���ߛ��7mrS��X��������;�+:�n���zz��;	�U����g {G� � ��%�з�f�>�6N��|�g�1D��rY�=�Ox��_-J�f|2n�d�`U��,9AW�m�ɢ8֞A���y�:��$�R�M9iw�u��y��tiӹb��{�UW�R�R�T�ݧ�@<Zvid������
��JA�=u���Y�|������\�gq�x֜��H�Z�3���`*^ڹ!W֪��z<��$�\Y�y�]�}�bC/S��>�\�ٲ���/9u�rTU�2�k�����H��K�V?��r�DW�<�DbH{�8�y���p�5�f���vg��$�o�^�Q$,=�G&m:C�R�G�@q�ތ���#X�F?�2vft��Ȓ3����\��可�pEhkWL(��Tg��mJ����ذ����y� ,��X��8�#��A�0�v߿�ͣp��-��K�|�R�	�T!Qi���������)�e��0�t�)��B#��L���iW��d�����$�_����5}�kq�}JK�?skz����8�KP�`"Vml�F�*̰�\8�T8[���쓆�@	5:���=�������+=ۙ�!�~�����U�ҕ[�~V�6��a�.����3%y	%y��F�TZ�L��I����f�}B��|SQ��#�����N�=gҗ��s���Ǜ�Qd4�r���J4��q����+�7����s��Z�
���=�ŗ�0��� V���5Z+j�t�y:��h����� �,��ƺ�ӿ��O��Q���ΝL�}��?�!��6B�d[k�f� Id7��T������	� 5����A��c/Ö�)�ڀ��fW#����ey'ML��[����s��U�w��8'��T�d�FuH�8�FZ�ox�yE�T�[��avS���pH��fR�0#�(_�F�yz�Z0[�s�KΟ71��s�9����<�?�)~��j�r����V����L��9i[aBmJ� W��9�K�9�7�H�Zrd���?��xN�k����{��y�V%$x�g���f����ؒ��(N��C�/$i��;��X���Ӽ
�	v��"[o��<9[���CV!(��QbX�c���F��'�f3ϫ3H�4�1S��o��P�K�Vh"VP7ZF�$M�fTvX�]B�L-�{�l�2q�2cb*� e�߉�I�_�*��6y8|US�3�2*uC@��{89V)x3`�=�ʁ|�4����8)�C1��Ř��9dJb�,V� �w�ڌ66�8���9���$��e�׫��lb����\��<s���
d��b��/lO�n���mJ4Pb�X~�ͱ��M��ϖ�G΅���:���ft��y�L����R��r4+ �!��J�׮M�����>�����J��z�^��	�Nte��!a�R�"K�E�rLDw�W%��z�jq�Wź��F]�ҡM��fI��<]1�!�t�T��S���J�P��3g�U��f���SN�u��WT���Ht�Yz��4N�Ĭ��eE�)�l�H����j�@��k�q9�C���}kB_/
�'��ʪk[�S�k�B��Qq$ˏ�����q<�Ǻ��L�&�})H�v9��g��>Ƚלw?��Z�3��}I�&Q!�,7��Y`ђ�|��������.���޶�������U�7%��m  ����:)�����t\�q����{�>}Z�%w*�q�������)gPw)�꒵�$�+mK��Y��'��	A��]@?Z	2;�NH���.C~�NQ���� `YV�����|�N��ڙI�Y�DLqs��Ž����$����l J6�Jڵ+i�A#���M氣Z�-QJ3�Cp�У�h�F�Vy!\;E[�����5:H�ݧ� ���.�E~5}�G�}i�J�ܧ��pg��9�)k�EE�
a�.�"n���x��&���lR�0!?�3�;�.�_o]��Ҳ2�>��E���cXdn|���>l{���6�͟��w�:��Թ��a��ӆ���sRI5j;��_��)E6�rI~�{}a���~x�*����`tZO���Ri��X��4�M���%2��|ff�^��bP0�I蛯���\�E�����6��PmfWJi (Z��p��:Q���M������3߮+Luܛ�5Kb�F�L�1��zg�]����5�x����`K�0u� ����k��/foEˌ�K�][�b2�s�3X��쐏��N�P�9<6�Z@���;>u.p]���@��2�R�N?>4���ϳ��|ij3HJt�1��K��Ċc�'��ej�v�x�)�8?m��ň=!F�m|����l�t��ycEy���LSs�v�q��:=�ũ�f���c����f3�X�He_�O��ҏ�!7W{��Ot����҃?��C�/+�_T:-}*�[s 2Ȯ�4�>X�?Q:����</g�����)H��NL�+��]⭜ҐѲ6��Я����\4w\zhR��סg�2-De2�KB�7 [b[Y��$t�j���K3�6��\q���h�� ����{���鈔f��7Q�@��=�b���`�i��s=s���R���o�)2�ú�����q��t��B�@�>��W������W50/�k���uC�nH�����ɥ��&�����g�����x��t���<7>3x���"qk�c���Oߍ�[i���ӥ���g�{�۟E�0�ǰW^I���Fsr�R��tM�W��?���j��zi�)e�x^���*K-ūf��v�Bd�ٓ��v�i��s��'4>�!�}s��8G	�ﯼs���"�OzY�H�����M]>zxqW-bj�ƚ]k����YOBmZ}#��X����@գ�e��]C�TvK�&a�'�ϒ"�:5+�5?�� ν+X�1����1_�ǩ����<#���+��8�U޿� ��fk��Zpq�q}�������w�QK��+�L���@�6V^=}�A;˛���\����+^_�N/���~�E}YXXh���|��%�ˡk\�O﯑Un�7E��xz�s�>_�j�dnU:o"\3��OCN2����|Y,hm��e��l�q����D}����B�����ڛ�K�ݴ��ݟ�0����LF��m]�[_,��?�qz�ߡ��23�&�*C�Jqj�n��1	���U�C����j 	݉E��и�T�!�����cҫ^�ҕF�JtTsV1�|��2��c��H�ҭi6w�'{���QuN�V%���x�k�&���y��TɊ�oLz��md����Q%t�S���qI���`�_�i]Bڌ�/��%�شΏp0Q7.!���y��½�T���A+�5u�@ ���l2��?��+��;�gi����x~�.��:���}}��w3/�YJ�{�-�U\�!c;*Y��ϴ�:��7*���,]{<���w�ӆ�]�r��/����}�r��EetS��ؐ�\"�ts��(w��[���*ʵ"�ｾ?�x�g��|�^���9��d���A������N�K��v#�ZLKK�pNN��|�{L�[�#L}���k>�nf��	�1��MRsy����B�q�C_�����3�|[�ɲ�#^�Z_��.�e�G��Ó��/L���{�=�T�	|��ic@�\&��{~l����p}&�847R��!����^B��ˀ�\��{;�j����Wǳ�Y�TA�ʓ
�Gټ
��=�~����<hC��o�Jrl4t�8����Gp�`0ɷ_��0�X�N�f�����^Jy�u�S��R��R;��{�!ۓt�����$���Zxfx��ާ'+���Ok|FZ���щ�=z�ݶX3ET��6|����?o�N*���D2D	~��n��[���4?�"�aN�z���KI�_+�|���mx{���wG>��K��;w���Z竤������Td
E�Bʟv�_�;�m�w��߫��*�{�MPj21���*��"*�`>J��k�I]ƃ��x=,��y4C�Kp���#Oxi�)ы5��K͔�\�B��Ev��JjJ)Bd�M�I�~��T�������A�.E���ˠݮ��U�� �?����qK�z�Ƚ�/��\�~�:G��Ę��z!��������d�{z��[��n�0��;␁��5�+;pt��|$gzq%ygs��L,��d\�����L����XP-��b4�o�8j�wo>���)U�p��+t���N������u���!����.��ㅧ.�[�������oy'�0\�����给��[7�ޱ����g�|������<�"w�5mB�O��\�����<��|8��?O]���$��p��F��W��CE��/�Գ*#"9W=[�..�0��
���2�b<���\t��sm��^���xҷ}�8���
�+�4���
�U1:g���+U���w���1���3}���A8���a7 q|��C-�$^���ӏ��.v�Rq�����+޳���{K���VA�(b5{�-O҅S5��m�g�- ~Ń�pA�� [�\��s����5kOݗ��:�B�x�_Z��X�Ѫٷ���;�%���]<�rpw����) �wc#ߟ���>vz�����f��������^�\(��]^,9�go��3TГ:$��␲�ƐQuv[���Qs��s�|גO��L��+�y��c�0i��ߒ��Q������/v�*E��@�~,x��&S>&�Z�?ty?�c���:��%#���T�T��}���RQ����&�;�o���ŕ��2��
x$��̊8�!�H��o�40F��q��BT��.�2A���(�r �x�׵�l�U}Hդ`b���]b�j�V]�̝��ۓ"���0���~=Oq����i�s�4@�
^�q��g���ƮQϝ�A)��WxI&�*+�HA���f���_�;����e5�X�����(<�q�]��~@u��c?2�<t��y؊8�~�e�RJDh{I)�,�+sy�,�*���ʲf~��5�'�[?�ܿ]f؟�/������fL�߀�[8�B�[���%��g�~��\4��o�x�!��sm��4���[��[��~[(���}ȇ�|�M>�H�����i]\�8O>U�s|n��):��C��'��G.��V�<I)b^��uv<�>Kk9����а�qr�(g��g7��j����s��G>��ϝ{���k>��������R�?��}��;d���p�L���RJu�h>y��k��O{�xJ� �G[���e�
R�K��\à����n]^e��3�pW����s_�9�}��P�Չᦢ�,�����A/2>�;��i)ڏx�H�ꢆ4
����f�W�T%&M7s��G���`�����q{b��!k`�����@��@fc�佀h�߇C�w����{/627Ȟ辤�ͧ��25�*������OÃُw��>6�
G�n�_�1[H��v�]�X*���t�/�U���CZF.M*���r���J���=j��o����O��jE��g@.\_��-kf�'��?���,����%�ŧ�H��'PjQK��ܮ�����}�Q§���P l��Z���o��0���J(1������o͓O�gD�gH74?�U[{T|�z���s�h���[����A}�zI����η��v[��J��~�c���ݔ_b��n^��k���[��l}<3Q��c�x�͔��V�)x^�go$]�c�3�ꃌ��#u-eHU��b��ɯ�F�m_:�k$��ld��8]d����8qh��d���\��?�
QF׭i�e�V�^$1A$9�I��;@�gO����\������\o���	j�D0�K����A��K	����ɵj<E� ��ׇ}�6������K�>�f$.�>�n���&Df���f�Ϛ_�s*	��r��J��߿C�j�Sj2\��~ys�qgG3����v�6k��������1l�������aܥ��C�u�Nw���4��պN�K�b=�p�lFj����=�8�����a�k�F�Ov��Ɛ����&E�.�ʌZ�>}�������?�������L|���%o����Υ���K%�:v�ϴ��~B?�g��{��Έ~��ӧ?��]��qx������i���#ж�.�P>�Oٻ���~nErOI%ߊ��~5�j�m� �}�ђ8ˊ�h�Jk8q]GbëG���J��Ёqz�Z"&3�u�_8�,˹�r'R+�s�\���\���Z�j� ��%��Œ�]�Z��<� �y
���i��[ kb�w������)3:�=��_X��Ƣ=��Ƶk8'���&Y�|���gi"�*¶D�<��MT�α��r��m�4$ً�����,��{�>)+a�|m����I��Mk���[�wN:�Υ���nÕ����Z}��w������wo�,�6��g�ץKcB��+�;��>��䗯�(<u���+Ŧ���+��ĥ�@�#Af��������s^<�'��W]�����_���}�د���Bf���/�9�`8��D|g����mj`�=�M�^��ѵ.��o�=R�~}��!N/��O�fq�ċ�w��'{�p� ���D��kfBƩ��&�5�"$�){���⠶�֤O�ɽOE�wf����%t��Z0�>�دف����0g��t���7���aq{q��R7���<]�֘|>q��І��f�|�ݬǕ��TX����͚W'��f�ɪ�J��4��j��ua�{�d"�/���v�L!�w-C�6�
�(��V���m��ę
�1���/V?�����:d�=��'U�L�4t�|t}���#;�̏��ʅ��| d������.�\c#��>����pvF4*WY��ʄ�<�c�z�����eWPJIw|7�|��
�aw�o�ɯZ�Cep��ߕҵ�}��vLwl�~���2�!|�p����I��6+]��������iUS�߃�K�e@��|����d��<R�|���iJ�G&%X�ws�lDA�{���M{�ϾƼ�?�StJ���J��o�9��X2o��l���{9�ِ��D��kS.&�~��se�Ƣ��!�&2� ��R��e�*w���J*��6G,�C�6��P��=k���2��qX��^ԏ9�G>���r)�w�3�pyO@�����Y=Կv�#���n�o�Q#�
�ZX���צ�Z�u-�4k������V[o��A��H�vƵ�.�?�IM_�z-����M�Y�z�2�	���|#�i�f�%FP��k�XZ^D���?�Q1"�zKƍ�kB;�����\>t���?�k[�.�(�7s��D{^Xl�����Ç��nY�V������N$�d�F�uw%\�{�Sb��"�g�Ti��(8�VU�5�1?;��FS�+�ktŃW֥��F����9&�ϡPc�4zbpQ�=���j./�q+�OǮ�����Y����7xiY��c0�b���ӹZro�&ո�T�ߣ[���DL�N�Aۘ��5�ZK]���tk��)-�����y}�is�Z��nKw������[Y�����ɻ�ϏH�_��z�U����#�%��i�k��V�
cV�N=?q�V����n�e��o�k����͂��7ջu�H"D��b�#E	����#��U�l���ݖA���^θa��+L���ܣ�yd�i}���`{4Sr�k�xB]8�l���JeF�KW����C6�֕	�.-�W�����7u�d^6	~��h�&��( R�}��K�P���榑��.�rM�z�Y����E��N�ș�?��~#Y���,�N�RP#�rFu��.]�=�\2O8KzFf��pKs���q.}.t�[��B"��e�o�~Z)L�{�A|�������}�n��0T�'Ap=q��cp�a����'�j�-���K��9j�6'�~6��ʞ�p{--6zC�Վ�����������hőT��{���0���6����FI��&�'�M��h�ѡ^fY�\H'|��b>cU^Y9c:d�����ݓ��~h�ډ�6�'E�w]\>�ǔ�<y�	�E���nz�BQ�~w2X�daՈBA W;M�a-��=�f�����Y�9��ÜqE���RG���@�z��g��X��g^���ף޲ԥ�*���XEܻ�-�G�����yU���U+Ѽ���Ӌ	����獸���u�n�
�A�*6��+~v�"K92�����M��{%<��ʤ>���Ėud�r*�s����M	��s��U��yr�;O�hf��V�CF��ZT�������]�z���JP�C ��c+�>� [��s��'��E�m�G�P�6��7ׄv�.r̈�pm-g�{�D�$����BTKK���Y@ӗ*�ةl'
��nI��6�f���� ���?7�k���ŸC`$r`w�����Pq��AN���'��MV�ci!�J��vd5.���7�@T����z�������NP�yX��f�,����2H?|@z�w �����0	���"z_�Nh�.��rw����+�bmM�����.��ܠ��x�ŭ�F1dI�nlސr�o}pLu�յI��97
�R�J?$���Apb`w��F,����Z#i��7[6�.L�bYi�`�/��h7�ވ:#�ךYD)%\��+�ƍ�Qs�[�`j�p��+�!u(�<~^U��1oc0̗��À��b[YP�3�x(��=C�jl8sՈ;4��� ꧙�!��X�D|��C�w֖hm�V�x��yF�א�UG��+�e����H�5���X��XZ~+�_�L��)L��W�&C��bKK���(ztHx��++~,����d�g�c3
���r���j
�	�_(�p�;%���M��9d� ��6x"h���?������T�R�%/U}���	w-[�9ܬX����}�>�&kO�����qf�wo��B��vfN�E�&k�%��Vf�� i8s��$&�^1�Rl���N-"~\��I���9����YF0�wL��S7�l�̦#�R[
z��焭����{N:�9��
�)3�ʴAa>�RW:Z����=�&o]@�
ˡ5w�2{�J����5	�ץz��Ld�u�Y����?�?g^�H�J�2��4�"�j�I�]R�ǰc�P�nZg{^̝>I�, �$;(�~s~���ޥ�޺�C����Q��
�n>��uB��&�C��R�4F�ME�>��pT�����ˇ���֏n{��N,K����yi�*/�pR�#��Y��+NeOS���ǌO��D������� �zb|�3��߅�^�T0[��O:���ӑ���,�Z$r�v��F1)�%9ːYb�᳌࠰vHPL>Z2������Zx����Hូ9� 5���[�}��(Vw!iT@��ӣA�>�q�Lb7�d\.�j�l�l]�� t��m�X�c/foI���S��G���]�͊�Mo� :ۖH&\t����c��F��s����Lݓ+Vv���w���`����#=cL4�bL��t����G2��� �:Ju��I����~��`�j�m����3�W�iRRn)y��'���̚v�l�=ʞȃ���q�<�m�3<^�=n �w|����:h¿NiI:7�x���*�}A�e��po]�e�R�z�R1�Aܖ8��	�q--]1��F[<��I����q����ڪ+!��Q(�Kh�'�A�9ͣ��_���"�L+��@��ڧ�7��Y=�]���+�����¨������
�!�Q�� �J@�}���L����P��QN���s�}m�*�%j�)�ν��]�k>���H��T#�;���v��� i|�-�!c��U[:߉���>�5��/C�<O�����=ϩv��!Z�Ǵ�0iXpQBU�W�'x����=�ߢ�E��b�7o���3ԍ���!�	�$�˜�<~")_DώA�e�=/���Y-�L�P�\a~�N�)͒Nd�?����ռ���1>����S��P����]>�2[H��c�?��p��*R�+��Ej^��q�M��8K(���E�א�-��6�����o���r����\��Y�%��"@�6�����=b ;��,Dpo�(��{.�]�H����������i�0����Z�};�n��c���n,8Y��n�3�x�g!�$�>`l�KY��	�JO#3�<o q�6��Ob]��)�<K�Ũ��U]�R�T��������ط�G�}v�"��8�!�J"&�3ɺ�
��b�i/��l�A.��f���zN��l�P<�6�M^�F ?�0�TF*���h|��"ؒX��kY����W`,,.�jlQ*&�&
�����wF�K[��>V�	1Y�������9���]��i���Lt�qI����na�Ť#�h�*_�A�W^x(��B�b�7��Ϟ�*!q�<B��і�"�Ckh�8��^��a1�>�(��VqA 6��p��-��|��Z�m��	?)�����j
�a��%*�&� ��;�B�
��H�d
� 0L�P�����s���4T�'���?��Q�0����rZ���!$�O����G���:�pk��[������w��J�O�O�㐿;�{��= v�S
�s��Zؕ�i���z�?�t?G�(67��3�.��
�:������ZCu�[,ۜk~�A~����u��.2#ݺ�l�N����R�6�I?5���ݭ�8y�/RlM�+s�tg�>�Q-�:��m����k�70���_حݫ��
�G���K�W��~�Z�Qga���!GJl�2 m*D)P�ʩ�L�z�=�}�����9I���􎂟6���V���d�M�SL�Q���DR��pz~_��B�\L�0A�!�ղ,}�=��-=�]|�y3��b�_"�}3mx�XB6���Jg�Pj�Ux8+m^�\W�{��:���|��R�3�W�uS��|9��\�U�¼��ұ�qY�]S��vQF�#�&w�-:H!�}o�.���4ʆ8��Z+܎�UX�D`�¡��:��{��-�sZ�9U�mz���(Ѻ��5 (���l@��S��XC��I311���ro�[�w��N����Vĝ�|秷��T"Y?,cx�� \��}(L����C¿gVegY�س�v��<�8��W�f��	��_���2�s�GDP�o>��&{Ej?����!go�c<MhB\���!�5z�4dWZr�wt.���ŗV�^�ZQ�'Q��I��s� t&Bx��ë ���%�/ߋ��Rn��a���Y��M��[�p�0����qf�Y����Z�]�m@�v�lHm�KU�t� ZM��U^j�(��,H3|1y3(Q��
������w�F�q�B��'��Q=���=U@c&^���@���,2XGޛ�Z���w�as��>�����QWuQS���56�����f�[-סG�O��A��������jgsC�-e���W|<[:�`ݦ���	�\`�Ei��G���X_�F~�8�	`��V�.{>�����3��
��*�pt��P�U����_�[��D����)���N��ŚU���OΛ�.��L��n�$�R��{�T�	h�M^d�,�1�!��;GZ(h?m�������O}�/_O�m�q� �1A|�\�'���|�吵��%��(����<����X�Ө~��K���^�ձп/0j���y�1jZ�� �VYM��j20H�>{��@�q0}+ �JKŻ�&�-x����^1��8S؆;��5�Ԫ���OR08��mśK^SL���Q�\���������b�&I���p�釋�̓'6��M�B.?/
r ����3�J����d��O^+'�������z��9f�ۘ��M:F1�(	&y�&���V��Wj@C��5l��?�M��E!#�b��F�],1�Ƴ Y��.�|����+�b��Uo�����Bw��սF��~.��`���lnZ��M���x�qH���~�w������q��`촠���������n�����l@��3A�	�ʵw��P�D�V��؜����R��]�}?v0%\�j��o����]b���
x)!Sc�3"�����V�L���W�Cx��_WD��d�'�E���A�
C��kN+׹C)��vx��Vh���/���^���:��p�E^�8"���xzҗs�h=l���86��X+��4�FE��_�㘻��r�*r�;��D�I�ǐ�y�m� <p�pEp*�2��kWIx�Smu�k\`��Jb�j����3�F1!����<��nC�0����:OZ�ij��ߝiy� � �Ǆ)�P�0��ia��F���S��)c�-�4�1{q��A�� ����umn
j�aG�j�!K�)8����$�N�Ȍ���c(u��,Oq�r����h��G&�5|4d3���L�X��`H�W�L��^$K������F��R6���]C0���<;��	90 ��:����C�;m����/Ȕ��&����3����]����o�o:L�B=��}[l=����D�䇷�t˶���¥�$��1��/W�fT\]_�X?9���[���u���OvAJ�<�]ҫԍe���b@�rXΤ��g���\�/�Y���*��f��#`s�i>a��~�*2����V��l@ �x�/J+E�=�b�]?P�:��U��x������5+�TM�27,W柙�����ʬ� �X�؝�ۇ�C���T���F1�>�V��<Ħ��hVN�t(� �y&����f�(D���Jf\��)�]���)�I<�^��<�桺��Nzj�ɻ�%��gr>u����R��x�w�>D7RN1tY�tt��)��.B��_;�gK[ǺF����R�β�NƆ�7gwT�5��9K�g�W
N�r���"���_$'���գGjv�	��s�4���!`�"�q2ّ���e�t�d�k@^�����ck� ����AG#,>@�AI���E(������*Fy@aL"|�R8H���Uɱ�c�S�	�y}d)G��.. x�� �~e%�'K��_�؅�&`bǇ▲I��ө���H�q���e��%�&�
�i�c?��85���++�%���5j�]����h/�M�a��s���f8"��;����'��Đ @�_���iQg�3�~�5Q�hI��Br�6����kD�PQ�8.���̨���by~�J,-,b�(�-v�|{�v���rwZ�\,��X��b�K),���6ػ�](hE���8f&o���Y�N�k����ڍAӮA�4����o�Q�|v��gJCxM0ϳn���)� �,��8���(Y�� ב	����)>1�H���(?�[��\��Ӆ} 3�������%r �pV�tN��T�2z���h_���ݾ�IH�P"y�ZX= 3B���7ޏ�Y���$�������!�ւ:_'���{����W��j�[~�����p�7��z�/lO|��b!1V��2v��aE�EEi���W_W%��i�8�*�!�kd�=��ĺ}�|�=�]�|$�����Z��P�,,
���`	�]�[�7jV�"�9�����D����52�(�&X�3bf�d{.��¸)���nc��Z�:��t�6lZ���ƹv��XJ�󪢺���b��s=T�W%�)'�~������5Y�րn�j)сr�`6/��(��(��
���*;Z��=g��LLf�B��W�K��g [�G�ic*����U2�B��f�R��I�^��A��6J8?���r�ʵ^rQ	�oE��ڟ��/wN�1Z��;�.�~�>��^�{���Б�p��� c�Z��@�+'���`F���@��x=\�$�)��$f��.�T1���!��^�	������rL]Lawzވ�?x8�� 
툢�m����jt`�8�Ζ�t1Qw���XܙЊ!R��7��E'Cn��I�>�p�r�x>���Җz�/D��̳���M�v�-�e"-�����Q \$�1z��v�������}F���"�{��U��� l亖�[0���K3�*�%D�f��bLH�;� �����>����e!��q�JP���QG�*�ؕo�c5!^�� 8������3�����z�R��Q��*�3n�o�UFr�r{< Vح� w��Q������$�\�$�=
]�_p|���rfԪ�3n�wO����Gg[�"b+/��I�������p�������`��h��E!��!HP��q%�፸���1ި��O+�Iߝ �}��oC��	�����'q�,����w ��z�6�U\C���_�\`hJdPP�<Z���"�X�:k���<૜`-�|�'A)MxN&�}L2�uEç�)����w���Wi<k,/��>�T�9�^' ρ���c�iȑ��pИ��r��9ӫEj���Uf���j}�n�j��&�F�O��C}�1g���-f���)� �~�u�x�Zj�%M� �h���������J��w�2�ڶ&%�ห%��[#ʐ�Y>���{H�-�)����؏E�0x�؄8VS�5�_E���:��r��T 6�Nh�Mb�Ǒhr�k����qBO�x��Ћ٨��įz���h�T�����i��.e���P�t���f2�B}�D��+5hk��j{�� ���e�x�[�������@�Z�W�>�:���NY[��h���˟�=�y������ߒ��<�{�RFR7�j���H�ͬ�"�Ǖ��/���x٭�!��$�TqC{�|�G�S�)Z��ߞ�S�+ݾw����ƙS�Ë��E�:+��>�&/��l��t3�@[EU۝v�M��(II��^�JC��o&d%u���ɻ��>r�Cl�N@����;qwa����W�
TdY�E^���z�����V�#v����Q|3�juJjfa�[rQ�4�ĹI0��f,=S*ǚO8�<Ep;�����I7��iX'N����y@i�\C��{�T��X*қ ��)����E��a˞�t�tjX���̷���D~��lق%�� �-�wE�Ͻ�3Iq�-ݳ��Gmv�t��iwͬ1�����A��W+�� 6(�N�~��8�q.���d�۫��y�j$z�3	O-��i�=�~]�Ը�U�%e� )�{�J�� %��h�@gKKK��m��Cs��Ga��A�������T�+V�O�����W�I�����A_�|p�Tu�V7��؏�G0ٹ���
�0��>���|^{����XzzS;I�� h�yY�y�N�\�.�1�<l����S%��q�ÄC����vİ��P��b!tu3c����<�Q�ȗ�C��Q��z��IG��%G�+
Zz�����](�i��er�������0�ܶ<�Wl�.���`뼳Ԍt���&6!k&vs8�C�C����~�S�q]�Y��Hʌ�%vRc*�}P�8�d�����A��SE!��������.k:��9�>͋�����������C�B�ѵD��-�R	X���7�m�?�O����W�xZ$N����g���R/b]Qէ�"�)�g���r;ۼ�Ip�;�4a/���?)G�t�Ũ�V��(�?BPF�O	V���T�J�Դ�<�6C��g����r� m��f����6����K���	�������fK����f 5X���Z�����O��uC\�7�Ry�K	�4Jڨi�3�߳���Eh���^I��i���)tP��u��qn��M�/������:�yH�/�o���/F�u�a
��T{�g�Wd�L�m�4���Κ꬀S�a!��z³(��"��bk��I�s$-��fYX� �WJ�]��ܢq�MXP#�t���b]=����,�[�BӶ�V����1�	���LcB���6b�hI^U�o���m���r�X��Y�v��'v�)%��Ag?"��p�e>��9��h�a)��(�8ϬN���Yѕ^h�z���{ ��V��� 	J�'m��-6��7�KH��@!L����C�P�C�k�3�"�rY��Y,ځ�*�G������`]�F8_x��a�4�ߩ�_��~���"��	���%3ǽQ�ಪĽ���T3a�l�Y�]�;IͮH;k28.�����\o|�l����r�c���x�P�������u����zs��f�g+p�Y���I>���tu�o7�ߏ�v��6�c@��xΏ��4� ���5?޶�A�8�LG��z����/�|!.��%æzx=o�aKqЊR��S[p��Q�n��N�P�5>C�[^��>b �I�^	���;��oo 3 ���uB�$�c��̇�ݢ���SXq��3c\$��)Pq���!�5 �c�ň�����[��݋��w
f���S�������^'�����"S ��7Vս��}�T�Y��=p�!(���!���=�tr���H�X�M���!F<ZrV^zL�(�1�!(͈	z��.[���ae�Ưg4)7�����u [r��bdb%�I����7"���vJэ��U}_�Q�!�����5�XQ4)�D�Od趃	HM��	� ��ݝ島E�7�#��j
�P�E��9a�V�W
�'��
|T���$-[t�������ǿJ�n^�թ�ȩ�4S���̖R�#�i-�~�^	U+�Z�,E�ڿ�[obJ7��93����D8+��r��%73NXP�n�?kd�6��<zlWI�!�[A1�I1�\�Ńb��J����}֞�H�p��	�
921x�{����DN�Yi�R@T��3v���LA*���rQd�T������p�7�$,gs�Q?��yO�&���ю�'G��u��z��]��8�R�
Dl�ҕ�?Y��z�2�d
�<R���4$>�5(e��0�%�2�5���C����g�A��8�[���!��
�8�cV{����qY}��N×�D�a��<"�/�9�L��l5���Ҥ,����~؅��0�m���4s������W?W��}��w����ųϿ=�y:w5x��Ott���+-����~|���C����#'R�%��ѣ`�+:�j~V"0����:�m�/�=~
Ͷ4�|�7z��@��~5Ww#&Ɨn7$&�"�%�-��J�q� ,�yp`�5���Mj���57�?z4n*���b�@s��4!Ȯ�V�j�J�r�㪴 �;U���>ׇ��	]���suv*�F�L%�h�\8Z����se��q�)b
7K�f��_��;�{u�}c����wPA�s��)��t�m�x�����'�+?�.��]!B��YV��.G�����FMQ�te"$Ϲ��[$�2�e?����[�n�4��<�/�IYR��f��7���xi����B!����l�
]�N�'�'xY|6^F���[��*<��CbĹ2�}��X�/%���v5��k-��k_\� :�P�˔�(J>M��B,�q1Z�{ɓ�gJ^�g.
�D��%��0��N�>F�/6������� �5�F�2U���6Ǟ�~���Q��7�_�sr�Οc�R}m���������r�ʜ�e���F�.���A��I��Hɰ�W�x]�zM_��U�>F`���L����݇�(=��rz�۞Uz����f��1M[3�S�.����f��d��t�K�u��߰�Eصq�#
�E�n�����؜�d���kzM��6g���*�|p�_�-ͨ���k�-�\e
��ìv�֕��̧�r�<^ ���O��;�tys�p4���Jkֱ�j`��'v ��;v�;0�o8r3��b�}�<e+�?	�]O`L/v�ONN����3h~���aa�	·�f?{;���'�u�W���劎�hqŕ�a�7����1@������I��W��f����ؤ.�Q,{�*��c���'��PM�o�`�C����+�!�t��K�V�_��*�i<r�W�rP��7�
1����:�Ң�n��Ȼ �{��[Toǎ�J�t]gH�������U���l2��K�� �V�s~��M�@��*�|�Aه��"�� �j�� ��ϊIzW�ƻ\�E�I4�0صޢ���R�˕So��y���$�D$Ze�ɷ*FR�~����Hp�nRL�3c�ⳅD2�ys�w�HX�^�T.��bok2����V"3�W��!�N}�i��>���]�)Z;�Ҡ�օ��.��̜b��p�'i����/�m���ɴ�,����;����iu�m�I�A�ʓ�?߆�kM�v����j>�:h����F7�0M.;��>�I���7���6\��Ƚ�������?l��?�F;p+ǂ#�$�W��rP���Z;|���$)�����Tm���;�BĿ'���Z'��n�N�_/�!3%�|��-~Q������y>0���|v�	�(U�E�y�G=���U�r%���S�'�Rc��Wwl�w'��*��Z`���\�Ӿ1�>e���
�����f���z�.���!�uߩ^ey�g���<����Ha�g<@s׵�۲�=q�Wo�+��=!jc��
��ҿx����7���vۢ���gO�����DDC�������8�~X�1����]��n��CT���{�;�}	���~^_�!	x"��B����.P�ԧR�%����qr�Q̺�.�r�� �R;�����.5�c�NER\���4&Rd����V�i�:����8��2�OY�o�!�u�!���s��W�k�7b�u��5l���/���H{��R�>�'���lgG�[VT%�n���hzW�̌1��*bs���ԁ�`4?��g^=�8�س�|�c�P����'�~�����j��>D����e�	�0[3.�q܁B�~�O1��/����4����"�}�
�#��b�f5н�S�a%���.��b2��p�{�R�	� I5�QS�t�Ox]~k%j����yn~1�AN����������_���)�9\�̚�X�$N��l����h��X����4I樌���3&���$��68���_.DE`Ik���c��W-�q���H���&N����S�])]��`a���#����&�u%P�0�:�E[���x�.��[:k:s��D���n���������4ж���(��#5Xz�E^�X��������=8�m &�4�w��Z�3Mso �[����7Pu��2lu}�*we�\z�	֥sZ��؂��p'��p�@K��1�ݴ�i2�z7�j�UG�z�v�Rq�|���ѡ^"�AրG�HM����r+��[�WiV�����}���Ԥ�� �X�t��FS l���ʹ����ol����z�A�.I`)0P���Kb.��+�dD�W�`�p���J�=|�֧Ac&V�9FJ�P�$x}%
�"?�Nj*�s��ӫp�MGD}�\����)�/�2����s�P�qpMP��f'b
d�弫F.t6�l��#eЫ�s6ByW���/��D�B0��^H�ʖb��ɑ��y�QĜ��с�$���������0����!a�G�.b��l#�w.yo����\9I/��q��+MrA�5�G�|U޻�F�q`�9n�M�2�Q��~���@��W�J�`~_��G��B�/��u��m�"���~��K���ӕ8t0�׷� M�*��*�^b�D�+h
��%��WM��WQ�:�J�Ƌ�c��]��U��_���=���ȓ&`�8P���cu�m�!�H�R0�ȷۉ�A�Z9VDKO��,5��ג`0	΀������x�Y�m��ڢ(��,{9�ٖ0l�_�~���K&ȋ��7R��Q�=D3j�E��N�R��]�[���J`�r�R$4+=H����w�h?M=���W<�¨�\\H�����:H 7:�4lK�Pa1����a2݋�Tظ_�zKޭ}���K}�5��_�6p#WKc�.*~��<~��㗟N,���ݳN�Sڏw�������v�g�e�������¯����z������P�|��'	�:���'胎�Q+����Z&"��Rl���1�z`/N�E&_�8��	.a���F�[}4{nZ+�q0y&���w���RȨ��%�K�}���|%��Y6��1��:hh��<�eX�m�=<00t7HwH��twʀ�Hww �ݍ -C�JIwJ7����~�w�s�s�Zk�3Ҭ�	^E�?ӂ�LLy[X#n)��b�oL�9ΣѺ�P����S�$M�f'���x��F�wu�+���m7�f��Υ����H!e���Y��i����Q�/Q	�]察�G�Ϊ��䕵R�PW�WHƧ��a[ ���V��fܗ������}�-�~����S����'�ּ����n������+���aK0��\��턁'Nb�lS���m��������82��qB!O�ˠXNl��<0kcy��Jq=��0�2_j,CE�s)����VIP���k7�:�m��#�_8��:��7R��:R���v?.Yo�]�%A�)�ZA�sӒ k��X��V���-q,�B�XCe��� �~O�0Z�ۤ��!|�5#}෎ě���4�TI3�h�4��>GT0��s�6z'D���}C��K��U
�(����E���ym�7B~���g,��g�N�иa�T&���:V["<|<l�|�Ҫ���^����-n4�?�9T��oZ��m^(�v"{�/;��~Jx�]S�~�����m.ͱ�;�"l�&��f[㲊!I�iK���!�������H��A��~z`�Ā�^Gi��`|c�w�0�{�(�3a�ڝ�Ԝr�p�D��r`w��XكR�X��[7
Q`F�t�e`*-k���<�SdeU��;�E��a�ɸy{ť�E���t���F�z�qnbc^>"e�=��[�Q�WV���<�W���Q��D������+��Q�}��fF��ze�)DG�J��rT�V
�gt��i��;%?�z��y��� uY�߼��S����?]k�8[��ImN�������>?�2�rtݚ��8����[9��V/OcJH3q<�)��z�Ѵl̺�=�,	l(x����I�����ˡ�C��	�y	.�����uiw��r@����{3��9��֕����g���.Yv7<7�*�֎WooVN�.�/�ST��l�-�y��iil���{�ì����E���@�y�ϰ�޲
��@�	'5��t8�����*�%�!��I��B2���'���~+�����7q�y��n�΄)iw/|���N��/���TE���|��h��-9"7�q5-5��'E��\+{��`q��H��͂A�735%�O`N�8����������t��p.g�/��6N/0o�-GS����V:��z��,{�5b�o�6A�%1M�0�2��[ݵ��Й�=��g*,�	Ë�Mص
�(9_ܷ�2՜̪:I���]�����H��z�o�~���p*��'B��%�O;X˃���v�WfßG���)WV�N�g�<���+/�#��c'-h�C�r/�C�7H�k7���>?���M�?8V��_*vd�<ך/��|*�د�X�G��%�^�x�ׯ_swK�c��ܜ���<�}ؚ�~v�<Ѫ�(D��	Η�ǩ���Y��@�lә��mʋ���0 �5@w��;C�fs\�0��,H�!������]ޭ��w��"��3O�Mh�r�Ƌ��4��0� �N��̥:��dI�~Q��7O{���L��ݺ�tϥ*N�� �[�<QJh��X�(��[�X;טA�<���b��ݍ0�V����У�9a~���.���9s�������+<V�Z�@�"v j���E�5�R�*`͒��!E�º�J��D��'ق�ajy���Q�M���@md�g\$)���v^���'�ï'fhx���밪����V����v�CY��ر�ޠCs��ѵH O�qڷej]�ݸ9�#�v<��h�����k����Ir�<�B�� Kǝk!gכ����˚J��ȇ5~'�?B�8�Xf��<T�#�f��.�w�-��{�(��~�}�:�n�C]�-���66H�'����VJ2�I���s��L�̧j�J���iw�$&��r޹쨉75��qX�z���𝦸4���5	���e�4�|&���>��vCb9k߉�ͱa��]�h�)��qJ�4�꡿yb��}#�TԳ�,�z�S�\��S�X�֭���]_F�8J�gOiU�.->�l�_��p	GP�9:�]��k�{A��w)����Y�!Z��J\~0�}I��ə���^W�B����Y�:�ӛ�x�[��*F�A�7p ��t�l�]b!�1�l>��k޻9/��P�O����O�fڕ߮C�,���oWo����([��\(��I	���:�|�wR{�����S��|Y���M�fa��iX�$]��eH��A���p����+���t;��K�S��|%�f��qu���N�dµ��!��di�Qvʓ�������ǌ�K%߅��aCvy�v�������H<�.^��=�o��%i��{ቚ�1bncؼP+��#������̺��o�C�W~�֝ԏ��	�x��1�c?I�#XmB��������c$z����vށ"؂�i~��:��,�sm�1��@[����u��2a�V�~�&���`�yD_|�U�[lYx���oBd~GH\�B�����j;�5���;��SY��*�d�'�h0Y���d�/�BC��S�����0�$3��f�_�T#���U����#�	�0�z���Үp�D������K��H,p��Qq�"θo9����D���lq�lD��7�"���3�w�&��Z������w�U�6�p;FY�>�9o[�|y��ilz�[�5S�㹎R�#_y-�и��:S��BjZ���;�0pi��^'\����v���b���%g%�I��}W��4�c�+�ؓ��D�RKH0P�	�k�l��$>�a�be2g�R�s�߷�q����ꉣ����?j�������!�5Yv�ca�@^�����O#N�����0tͧW��&�q4��L-/���|+�R�ͪ�i�H�9;O�?[m�c;Qi9�su�������LN�B�{�u�W��k=	7a ����3�h����{��n�����l�粳܅w����m�̦��Y��Qhcv��
��4ھ�h�z��~�aw�ӿ�}z#�8|K��J;co�w�w4'9p}r�S�V%������Gt�a�MTyHJ/vPhK/����'%K�Z��ʮ�N�+���xw�W8_t�C+�Պbt[��
�R�6����i���L� ^=����F~"5���E_��i�m?�-� �@[^�b*9� �$�����N�z"v�u
`����pFJd��&�6�C��������.����bT!���3`�|,�Yݹ����/]'�7+�/���/h�.���K'�7�[ׁV��j�o���\{��5B�ZAO�=Ơ��g��m�桢��'ʥW"a��y���uz����y�]�5���ai�4��۱~�����C��]�JՕ�64=b�g�j~��h���фo}b<-_��:�Ok^��-�}���V�ܣ�y�d��y����Q{��0��2�@h�����d?��w���,X湧܍��>?!?R�@i7#�(���J�'׮��zc�I]�\��n��C���t�&�E��U6��4�m�?�x��,x�ǌ*0>��\G��)�"[	w�b��Te�5W�����3�GP7�*�o��g�Ӆ����W���G"�7�*T�Y��&�NU��o���C��wmB%�hs�#�rC�HG�zl�T��p�
Z�Y���4-�ҥ���%�zz"N����)�Dr-���9\$�1�)���B��$�\��u��L���1$�n�f����)C�9��{v/?�:���w�=�mVb�S�%q�/Z�oZk'?���p����q�A�y�I̓����7P�9��o����Ë�
���O�Օ���ӕ�f��$����/GT�Z+�O��?�:�^;t�.y����9\�7<ˇ���hr��@������󭮻�*�f9)M���q
.����9�$��[��6�2�])H׀����0�8Ɠ����	҇vPe|w�(B/ n�.0=r�`"�>_�Er��I�
(E���2HFJ�4�%�
T�K4[���vo�w���*I�����Hg��>H60����Ϥ�Y���xz]f?5V��>�(i��|RDc��^@fRfS-���Jf�C��l$"3>�D�&�+��U?������R�?�M���I�̨K�ς��]ͣ��akmX��=v�{]�ׯ-E���A�^[B�~q�6��0t��O�8E��/;�w���B��Ϣ�k{+[ݻ�K��o�(OV��\�r�y���O����w��;�On�^���DQ�{<�>�ͬ9��^<������=����=w_sk�_:!���{:��kɡ�O�{��$���i�}g�����ɶ����kJ?~%_��^<�s(Z��߲5v���d1V�q�*'�/�v�'S�]:�6�?CbP�L�zlW�}�����G�����	������Y&6:���y�.�O��>Y�kx�0�Q:Y����bU7y{�<y�y%���-7�9rd�k��f��)9���j�x��rKV�j���jj��o52�|��ߚ�EJ��vq������\=L�Xh�����D��qµ�N�C���|R:/+`c$�"X�A�+ӂ��y8=NBP�5jV#�D�{ff+j
��5��ǁG�y
�� ��3+�HXԉ���6��X�������oyk��(6@y@X�O����`�YD�N��ќ�7}�:�;/2�!i%�נ�m6�b@)ɒ�m���_�ïԬ���J�.���X��������Y���[��Χ�� �i�	RY�i��F�I�%��c��ؾ��蓭CϬ�a^k���0O��aK�K�{dܸn-p�+����8x�i�c���n���q�(��3���S�d��%)ou%g��ӳ������?�}��!�P��i��!�}��X?43�6��I�wփv�h[�vtc��r_W@�Ԕ䬯R"�G�j�9��[����=��&�`�o_׏���[�oX@0w7PU�U��a�����4!�0I&jlk��(K��Uq��n��֓e�ۈf�2\9�&�U��V]#�XJ1Q=�0b:� Z���yw$��0��eW��&t.Y�h;���Mot��`}T�1�DxO��A�����u'E���� ���e�ke*pk��b.i쐩^սUb&m�`�
A�����x��X��u����2��[�m���I	fu ����%l�W}`�6r��Τ�\bM�0��B�6!��cұ�[.��:6佁��ި�tO�:E�(N�e��"W�aH�墤�*�:^����$���m>�0�0���!o�Ŗ�9�����"�3���Rڲ>���7�3Ұ�uO�򖰏�0�ֿqzC���W�
��gW�3�}f�g��_����s1Lq����*�2y���������������[4/.E���I�V\���az�}F���¾:7F��Ԑ�ce������V����_ⅿp��"%�֨=�0ޘ�ɀ��$�oV}��M =2��C .9�{x=x4�pb��o͉��]����A��L4�L8�	�.�m������g~f}�,��8I��,a	�(0R;��Z4 ��2��d���/���$��ZX� �
�ҵ��A�S3V0�+|����O�Q�a��dO�,Έt�ڢ���q��g� ����B��WH�������o@p��25�wf���ы.���!^`��Y��V��&�����+����s�֢J}�ɍh.�a�;"��t�� �����
K��z=q+�1>�.�5�G��{$Y>�<�F��ѕ���ͤ��*�r�y��H嗲��V����ѧүm��ϫ�c�:���� <����y�����"�}:��E�D3�S߹�/����Z����Ӥ�V���3ѫ4�\#(՘Nro{��8��V7q�����P�
��p��p�L1ˤ
K	���
�TBE���#O1.���Q+J߿aHVEK��!%�ˉ�"ĐruJpt��A����)d���T��*��I3�h�g4��]RĀ1[���h�^��/wc���'P�����
�&��Uk&�$ao��HE�^����N�\�>n�ɽ)�՝��{w�Qu#���nْ��0��J����� x=E.饟.͋`�a�ƭ�H�h���F�l�p�9"[qE����"_����p쩃�!����>O���~�e�_��,�Υ�r���3�UK�.|s��������BBW�H�����Ǝ���|���Ĵ��_� k�����&�V>���_�[��l�n���ࣦ���u����(	��Zc����ٱ�ټ&P�Ԅ�IʝY�j�+�yr����Z�@񿚔�#$����E�	�.S&�8A�K���;ݑcHE�������t�.\�[G��H���1�%��{�>�	$d~���ǡ[9����������3'��]G�M�L]E�]���4c���Y1�E���hP^��L����v1"��JQ"ۣ�^�p��s���(-@چ�덵M>�8=�XQ\��^�Qd&���,A1nY��$k�}S�?S�`��
��[㣍K��T�r�#Pdg�]E��&�@|� �N�a<K����*���_W��_�I���M��֍��Q��B͕Bg��g&�{帻���v�lstO +6F?�Н��~z�뛆kQ�,��]���ف��h�������R~eƌL������[���1Ob}H�"��c45���m�F�����-?��R���,����w��[�G�Kz�&�;<���}���	Nw���Nu�3� �9�9��q��3�$M޻�-����h��;4����o��o�+0�1��<�Ih>@��9v}ߛ�6Q���l׷B:��F��A�E��r��5�4��)�+����T���<ܶт��&Y!��)w]��x�Z�K?AJ��B�x��؁r�\�o�����{M8�Us���3`�!�G�E�������>j��j�y�!�݀���ё)\4򃵸�LԬ�E��C���l�eQU�-13D#�u5�˪B�FA��S蒤MQ�Mdt�<B�Z�4�G�^��M�{�v��D�zn�Db����m�%�A��?Lρ;.?ޤ���ad�ѳX��ƨM�|_�T�E[�x�9e7ʧ�78Z+�m���=�'�}��:^�1���Ĵ�k�37xRmE�hL��P�cxѪpx��S��z(5��7���V]!�Bp�@C��Z��Btނ|�f�)3"�j�1R���䯉�J ��2$�YDsn0���Ae,Qݯ�H�b��0�*ނ4c�&�*����A�q%q�r�H;ҟ#w=�0cL#@J���z��ɮ��!Hw����֛��t�G�j�����nR��ë��e�)�B�.q�ɝ�kW{�N;V�,��:�yWA�	���K�l&U�-J��{���2���;u��r3�����<a���#k��ۇ	j�.HQ������*_p����-t�0U�^�'�[p�]Q�=��Xz���O86�q^I=g:�;M?��������j��8���/��8r��c�S�1��tf8���4��x�P��5a���F��~T�
�L�'/�EM �Cm�أS�A��M�X��I^i��<�r�G�#��	�����H�NԱ�|Y��d��>�����W��2�?�O-�	�9sb\��O�t� ��`_�;.�2:�����y�܌�Ax<��z�w���|
��fsmg���q��Fz������0�	��RP���T�i��U5ӕ����0�������};6�w�^��I�ٰ���VVfR�4܍��t�`���+��Q��̔b�ߨ�'���d!BÀ�3ͫ�BͣT���MM'f��E1�ǚF��&U�z�e5oOI��Q�O������[jɻ�T!+�Ŧ�X2O)�WiG����S�7ɴ����[�}��#�ԁ��,o�g���ҍR
�$g�\||��~Ӓ�+i��yG�žz�� ��p�Wl��=���� (���B���k%Tx��P��Ʉ[��D�A��Ì&G�.�����>D���.�r/����*���"��!QŶ5�9�� ��~� 2h�/9^���hz'[��|�0��'���EO�[�{���3)4ȹ��?0����	&�u�Vռ�1�q��?�9�ּĺ��^7��F��|�X4E��l Q ��i�A��&j��6�5+�L{��� � %Cu�����׿_��[eY���q|P�U������(Mo/�
��(��:_�y�:�bp���&�h��9��e����r�瘝�h\čS������*�e��[~T�}�"骎EϝV�>\Ug1��%������E��Z��-��x2�oƻ��8��{�ԡ�.F�W��k?�	��a�a�8l��G����/�Y��y)w��2C�L/�z>@�D����߬q�M��q�?�Pڈ�Cy7����;�y��vNW��X�9�x���R�[�LG�8��A?�pB/���)���ɏ��&2���X�[��R�EX%`�H�𩒄k���[y`��c/.��5����u�3'?J_5F���^��U�os&���	ь󍨦E�m��=�w�(QK)$iHU�m\$TL2�neqg��V1��f2imS�u���5���X.]�f�pw��M�o�/j�Fp�H��W,J�r��C�K�gQQ-���M�R�7Teʊ�+���B�+I�O�+�)>d�5����߀t�,Nɮ��`|I8pW"�Wx+�ɘY��Q�q�W���V��(�5��%�䅷w�E���+m��n��Y(\�pq��T�h*�w=?Gό��0`Spp��A��zH��"U+�	p=QL�x�ߔAe>�`�2kO��q�WN��%åd�@
u���mS�o����Lg�����+�b���0������j���P� ���1DT@�?�#'\��8�I���Y��N�-�p}`�W�D�+UҘW��1���q<�"[ul3��G��S2���[U�^��T����DY�4%�� ��w��T��#|<�	_�*c�l�'K�dӱr�u0y6g�f�����\�a��
Q���89[�0�inI�#T�v������b\���s�o+������v�,N��I5� ��͢���d����9ӏ���"��)�i����O� ����#�9�2c�[�`{�=�j�������'A+�p<�p69�$����Cg�U8��G����I2�~�����7{�F���w�5S6�)�5��̾T��L�Ώ}|����h}��G�v��o��AS%E�V�]�;���7����@/@�l�!��[/8�R~w�2�I�_�!m /'3B�7�;x�>�������Q~���D+Gma�!zO�:PV��C���,1��ϡ�d��L����bxO&��a�
O���b�igI/���)����d5����=-zc�nh�������4��<�'���<4%	�.�YS7fU@������)M_is��3�k�4�M�t��2v}%$38��"-�Ga����&� z��E%w	��y�)��h �9��q�	��s(�A�x���������#��5M���{hs���q-ǲ���Pz�#H_�y���n���s�;qFp9֭�T@F����5m��q�1qer�*���O�^�J�@�8�V�}C2.�d6p~�P��� *uKꉏ�f��sXC(���$���������\�z�Ϸ�0�`C0km��B4����a(����dl�t�����R��L40�V��[/W�#�psjz�W�JVpU��3e҄f�ƹ� )�ه����s��q�;��9�c�l�VJ��;p��~��|W�9��ou����	��]gx���A�Z��j����[~�Au���&��CW�$�~e����/n�5��OO��5@o�'�1��0
����N��kE��2��@�-�W͠@4�x!Tp�O�&Z�0��u/�dE�c�������|�v�'�cT�-׉&p̏#R�� ��W�!��O$�����
e�����zӆ�#nc��X6�o��T��O��Qn�����^U`�Y�V{©g�0�W�nl�l�f�E{��Y���zN��U/�:���&Aw�\�|��,�J�"F���*��k�\��wJʷ��B��XMܔ>1����'2�7ˬ*�E����ID�}I.�ծVs���>�x$���F��g���
O�b���'�)L�,��\�!��CT8���^Q��9f������C40�x�(��������P�0'�}Q�-F�:bn�y6�����]x�Z�F.3�&A�[ȅ�B���<��k���fR�OV:	wd>B��  M-��BM�N��=��加b)Ξ ���H!͖����� �m�Jx�ku�hy}f�e���Ih���%j׎���_C]r���8W.Џ�2����_�m@v74uDU���-��نP�c�j��ʀ����O����"S!� ��P	b�1K�1�טw����a3B%3�$�+J����2�mعM� 	mk��g?:
�����*��C-M��[��
#��֧�=��b����4�ߧe��ʃ��P�cajlib��4��~N���vа��+$=B@���ws<�v���<M�Xn�Cp����P�!�>T79��� �X#. ^g���+z,����С��gҮ�0����8f��תN$���Fm)�q�&�f��W@��N�"�k��|�D0֚�(bM��f�2����1��;���U���D�����?��[�������@?�^�Ϳ-�"��	��;�
���S��g��CC��3Ƭ1��w�����L��i"�r7�B��5(�����g��`S�T揾���}R��1�2��_:�m_q(��m�U��)�/@�Q�xX��,���u[�pIQ+��?��Y{+l�ek'�q�e�����������A�y�H]�4VD�b�מ���N��"�7Rrp����`#�Y�֍���+�q\L.�)&���I֜�M}�2	�(��|h�:(�T�̬)�#o[��$�����_�p/%�=c|p�����tc�_Yj�qn���(߫�>��m�R� ��wX5��%�R�m�:DR��kϰ�@�6 �U��������B��^��B8X&
�D�-��m���E�= �㎭Ɂ��H�u��.F6B�
G�|��- >4(V�ES��u�zz�� ���lG �˻n�qCۿ��w`�&NA��?��b��H3�I@��t�ߏ7'+.�0�]0��O|8�
(�s=��L�a��}3H9fd�Mc�a�q��T8 �q�aR��_��: (��l\\�,�M6~�Ţ�%L��a�V)�B�I��H�P����G��\$�]���J*n��! ����@��Ə>5b�����'p�����`_���0¤B�&�V�_��*��Ш�R58�p5�ֵfY؈5�K?��b#\���S?��oH�T^[2Y�K[���6����N��/��o����K��L>|80e�=XEe���?#W��v c��"�hu�Q6X5��n͑�+O�
���p{��;����qVT��zb
���)M�9���Y���QxЁ{z�̸f-�#z�o+�EqLۺ���_<�t;ѺM�H��+h���ߦg�nn� �B�$|���U�8�p	����gա�{��7(M��w}ӌ<\˞�U�.r5�n̿ŅEw��UFCC��;�6��a$8��(��$���2��C��:.�v��rʬ&�Q%��nYB����)����3���}M�Z�3��͸���M\��qqSz��K�8�p����>~m:�`��w�vq�z-�=a*�����wֳ%�'s`RL&\R�N�C�_�|%�����lV��4@鲳��q�O� ���B�(�k��*�lݠ������"�?&a;2��[Ƕ�c�lRፉm�GɈ�;�0LS��D���"����R�ԝ, �d��'����HO3�æ��X�`O���9�",SW-b!��2w�h�y��q)&&nΉj�����n����a�4=�`ӫ��kl�H�!���8�����֨���Nq�|���=dG��>���;j����
�$E>����"�������v��rˍ�Z�'�2�_eO	�"{p虈r|o�2]!X����O3F��h/�z�`�;�ݭ�3�[��B����R��Mx��3��5qËѿ-�7��Y����2<�����lc0����|W`�Ze�4���M�W���K��|Ǥ�}||?s���w2��JW�`T��R[�?K7E%��6 ��e;��l(�3�͒5���l���r��r�w�t�tƴu�\ྜྷaM���@k�!�_�������H�F�w����(�����|��F���T����e�y'��۹�'V��܆���<�NH� D��8��6`�Zh��N��SXu iTa��+��C�����_9[���'\�]�s�
���i9m�0�K�Dq̓x�J�~�eR��P�(y�4��T2��3��!�WtWh/|$U���w��PY�� bn8.[?M�к8��1����&�[n��ߊ0̄���g��f��nd�g�iX/����<ýM������&\>�HD�"f��;<�i�k�W�hi}m�d����2*ŢtG6���e^��K�lkT!�#�|�g�1v���NKg�0�3ϋ���U�|f�YY"�N�(�y�{�����nW?����m?����Q:%2����"�ޜ��{E��z��^�7B��շ� *�g���Dņ���B�<q��يo�����~̈l?�c�2��2���ǟ����"�΅���0��ˍ}^m��ʼ�1�] ��������ArQ_8�0���D�Q�m(�Z#sk��	��o`��|��t.������s���w]?�Eۿ��$!pl�6T��?[�x��l��:֣�.���_�����?E��d��sط���m_�"pG}% L�Ąh�Ft�4�HA������`{�%��_�k�iF#ܚ��D2tp�^����L���
���f_5����#�[�"�;+���ғ�������%5�oK�SR5s����]z�E�8���3���������I�n�.�lo�k:�"�^[Iδ�H�z���o`rߎ�Nu��WW㿍W��·*���*C�!�X�p��`e��-��	^�<y"r<&%fHBetB�$��R��+�B1�E�����y��˧HH]n4�2ؗ3ZicuD�b6��4\���Q'�A'�'�*B�-�U��g��Y���h��CϮʏ=�p�X��{�_&"MO)*�; ��k�(����!"��[��6X�,��3͏�T=~7���LC�� x�R�����P��/ʯ�|H9���ֈA���}ϼAp�<��Y�ʕemPO?���ED>B�3POc��c�����"R~A�ӈ32��㏬(-�h����N����<j?Q�p\Bb�Gё%��m�L��_�w�$�'`u�&�'��ͤ���-���	��0Thm?A�*�*�"���po�0��*�W��$��%�#,�V*�M��;�Z��Կ&Oq��,eèǱ8.Λ)=2�gu7t�O�\K?�!�\�U��Jw��1ls�Vx^��	�d��Ðd��p�~1����B1��܀}օ+b�`� �'~�j�}�p�����>���l5eX˹���PBD�E�"�!��r�(��"ݶk�쐤T2��D�hI��x%t6n/�n��}x��+8[,�o���H�k��1���U�
����_�nrN����BP��|�>C���B�g����,�,'v�����r�uw����T��7��cSB=TU1 ��&y�z�P�E��b��?1j�̘�͖���a�Y���S�ʂ�y���;�A�J�����v���E��|6���
3Y`,����Y���1�_U}�	���8����B��9���{뉼Ծ��jyL������E�݂�b�nM*c��L�K)L���O�	yh!���ìy�`7A�h=t�k �(�i��M�?���^���<o���W��D��?��Wn����#ʀۂ������?"}�G��e�s.��OY�	6#ϓ��һ�dQ.Lxp�]5Wd_D��h���!��+��l���y��G�Zݹ�P��CeOW"�?�,f.�KC�w�XV\(�d��d�FL� ��������E�� �.��n��1O�/+=�\�*���P����>oȝM�x�,�ɱ����?ć����ѩ`ÁI�?kk�r()#8�|S�e���Hb��v�Y�Syvul �Y܍#T$�Yy�<��bHɜ�(�$�����CO��$�0��Ğc�qb�}0���/��`�"DaM�74����nc���1�����z��)�Y\o9B�O�A���N��%Eu��ҍ��T�<�{N�v�qE@<��}�~�5�������S�S��*G-J��KJ �u��l�?��8�Nf,Gx�Nr�F��v��N?�ޥ��K��룅1��jN�u�y�]� �{0��&._VXWD|�\�]�e�/[3E�>>��޶�]�%�6	� ��`��ҝ���h7��ҽHo̖�ɡ�*��R��D�F��%z�� ��� ?;	_����g?8#�tm�rN�Ynk����{#/f�~S�;��6{)�OJ�H�k֍�w�}�Ν��6M�a���xF�KI���د�4�95���E���1B�/Ncٿ֍�ڐR�|4�?ʩ��6Z��}�K<��ִ���h튑>�`!��V�*2����E���U�	��)S�R~�5�7��}?gޗAIK�?r���g��dЗ���z��j��l|a��i1���r+&�'�}/���վ�vԖ��>=#��<�C�	*��n`hخ݊皿��0Z���~�)�ګ%��q��#�?-� �X�J��^����I�i6W����X���e��G��q���8߭�|�3쒢�9�[�Ҝ1q=�6���o`$q)�W_�Sr�w]q��BrN��b�2h�8 m�:"��*�
�K�)0����I9,[��=�i�Lp���w�������&	��l]Ew];�[�`�`H�h �x���_Pڋ<F+Z Ia�����׌�b?�9��a�v>��37g���Yr_9T���6�e,�.�5��� A�?W�zViT�%v�2��R0squ'gk���b���!-�e��xk4uiE��3�$+ko�!ubGOΛ�Œ��ae�j�GӀ����eb��@Hw� ��2��d�i��1!���\��aˤȷ��1��#�,5;zz�o����V}��j������T���@�Ё�9`�x�}p���H=���Cp��h@54����^�B����7(��2���ݿ�(�o�1���?�e[�o?��(�(��xج[[y������E���􋄻8p[���x�&@<(���(C8��#�Fm��P�L�0���O�oV�&��M}�I��7��}z%��}}�.ϑ�O�I7��!k��{<�D�e3�l�I���������6zz4��y����vK;��A\]��
����#9E�mQ+);�'V���]p�"�h�<��Z�1ʶF���B{V��/6�v�T�������6����zń������)MWs�
Oc���O�tNM��'�ݤ�dځ����<�\�����$�d�,:�K�k�q�|��O��딛��ż1C�=��&�L����&J�'����Q���u��W�[�%��j5�*��+���Α@��g�xG^�j	�R�#hid�Q [�>�C�?�r�.���g���>��mz�v\�bYǉSQpށ�O���z��=,8�G`���;a�㝭2�`H�S5LK!����?���	#���r�3L����h����.H�^X�M�LR����h���Ɣ
O(�S���K3��'��*��D\����&U�E��E��>����v.��]��Zt���I�-�Bh�@97�T�����$�[��!���N��>�>E6Yg1���JW�!J�J�G}B���''
��n�0��'��8�0�;�r�8�0�:�`u���A����aZ���-^��!���4ҷ��7���qUG�ZxB����ԯ�}�l��-p�)�zN ���l�W>E�xo���?s?6<�������e�X�f�~���%��DcT��r�KJN�ɯ���-���{�y��>��0�Q� �9��`��5̈�t�7�4���NT�'w� 9F�Ùʴ�����I=�A˲�}A^!!,�lK����Ik�E�8��������X��|��<��=�L�
u� ����}�"����Li�Nq��x<*���¼��+<�<���o�N%!��G�O��a�u�WRs���!Z�)�>��7�<e�y���*e�Ѡ�����r���!���z蔒n))iDi�R��c(E��	�i�����e�=��<���־��ӣ-D��)�qd�����^��'��'t��E�&nbx���i(�H��`��aU�}���)�M�������[�D/�ʵ���7:uif	n�+|�jt����!%�)Ww������n ��l�@��X<�uG�����n���������ܦ�*p�a~����LF����u&=;�rWS�&e�7v�t���yH/�8s� �
<�C����8��z�q.\c������l�8�b}6��`,� !���SY$�����`S4�?L�c����r��rPao�BY��߹�^�(��)���	�<����:Ҭ���A'� %���Ñ�b�eL&���������5H(� ��J��3�x����l�ƒ�@�`��L=gͼr��5mGq�n`����L�Q��i���OVL��Af1n/W�A��e,�\�Z%F���/��vI��[J�Vv��
?��?���넒�"-�F���{���mF$Y�
���`�+�$q�慝�[�D��u�I�ć�$��)0$i��]�&�·ݸt?��Ѵ"������Ru�l)�ӗ6}���ϰ�ι���#4���M�3��<s�3�]�aב�D�E��/�U�S�����I��f�[���h٫iuR'�YwҨήl������U�y^©��v��1��nC����8��j��oxT&��`3��D�E5c"K�޼^���"�I��-�����;��A�g-�;���jW�����4��f�J�&Jɶ�J)���+b��F�MC�����vI@��c��<K�a�QC F� �=J�(?�o\A��e�{�\m晍��i�kjT��%�c����zc���h"�Uq?�,�О�+AyD_ER���x�VCN~���t(�Gg1vf@N�:}���=(�=�$��I/��*,A���S�es�Կ*�I-�ɇ�i�a�⵳�2�c(Y�zY̑�J>v��0�hgu���W�A�����`z5WA��ӻ��5��#�y�5+��l\����w�	���s��ǲ�;o]�'kL��
���Ǆ�٬���z�b�h����y~~ˠs����l��������޽N�ǏeE	�WP���%���N���Imť+b�U�,4��^��Ԣܽ�_�鼅S�>S�l*u�ĥ��މ���e�}�9�|�˿�A�|u(��U[���%�1�wA�C��_5]2c"�3��~ID�EDL���gaQ�'���@�{WH�T�H`'nw�����r�]s���gݳެZd�Y��'>�I?�]S��ĵ��J�LѠ*�L~f��W�\-#(�ھ>�2A���-���jH�������F�Mg���p]ie��t���P��	�e?��;�Kꩴ,X�{�	���CzQ�޾?�O*~E-�U�ي��ɒ�i1ne$M)Vl��ĝ�\#^��\#<v��Y��_���a�`ק�[��u�Z{�,X�������at���Uc-�^�wO�g�����toW:1��^<��G�0���1PpV7FyҸHRn�T�=����|��ɛ2U�qa�kL|a]:�w⪿�9��T6���v�M��Fv��F���՝��s)N��8��y�H�����ܧ��n�����O��l�Q,u� ��赲��]UO�|ٻㄷ]��J�AR�ﯷ2���0G��s����.Kf�󫺋�����T�k�_�EL��?��Ӕ��}�x���ƽE�����W<2�3�C�WO�:�:�8$w��U�����w�t*����h�����^j;*L�.��RE�ك���znr�iNZP�@M����
���,S�bM�,"�{�9W`Ti���%�a+��_r��Սgq��\��k$&���\��c��	��\�I�Y '��ӗ=6kM��ڪ$��ANz��4��6������i������xT�] �q��Ȳ�>�܂��D�����GQ��Q�6cq,Y�*�{���i��*�nᥦ�z��ɍ�/Zq��ފXy>k�0�4n��l�Z�Iڈ���&뼓���**I�r@�ԙ.��C�����,�Y�k��h�#^��(�W]eOM��T��Hk��Y�
89DE���7��0�K�j�3�/};�A�����<��k$����g$?��t���@+V��[w\�@l�l�X<7Œ���a��:7��"���z���#��T2������c�whᯉ�(�EU�s�p�8'?+��!�1�_	b�^O�6���=�i�e]KES�^���%ݔ�tcq��%&��D����"�P�A�>������9�k
�!�rl��Z۷�A��=�B�����-�2qg�W�t��-�R,�t���#�R�+
�.��팇ەG����g��H-Ɣ�uݝ&�俯>
F�0|���ol&�IQ���{)>/ݪ^D�@��Ā2�x�O�^�߻�!}MU�o$��DB���4�J_�N�sK��,)�ț2n{ʹlI�֧V-�-/�N��!���Y�9��Qu�C�<Zm*���-ޙL�bu2' 0�{kz���m�Ʉ��{���Ԍ�\�xU���3�Ք���a�A�j[*K�v�I_��L7�
�
�b�t��t"�!74��oRW����/QQ���B ��e1�|�m9:��w����0�c%���<��nM|�-��{��w��Эt����%��#��Ubۯ��	������W�|���b0M�M�E[u�&�d1�.|A�5��>yK�J;�~�O\��2
�B����|׃���N�B��H.����ɠC������jo	�3$�ρ8M�q��ڶ'��o�̦�d�hȱ��.�+lb� ����~4��H���R�uIci�~���&���X	�v���&ϩ�*Y�~d��+�S1�rVS�� �#xZ�l���SH%��j�?%��e��'����w"o�Z�2���J^t��^7�c>�VS8�@T��N2�t�8�}H0`����������]�֩�gF �Y���ר\}�Ab u	~T�Aw�Pւ�������e?\�����[)1Cŧ���̓�k����g2#�^4��� 㼆m;�`�Q�c�M���R������^8�U�JIm�HkC��O���O?�X�R������R�,�q�Hix_.����^:Y��������b���ts����w���s�Nx�;�2�	vQ�#���,!����*w���kw����f@N}���7�����7��̮�K��̴DשҴfPan�f�á4�L��ڗU0�w�Mu��{��L�rf���.*Ze�fk����O�����͔�
�HS��=�M����	MiԊTt6��$��~aηTRGk�����0���85=�}�Ƿ��%�o� �Á|��:�ޑ����GZ���?Ŏ�&p�MCI����hW��<d�D��V����l�'��{��>���S$�@R+@}�񍅜����J(���K�j�S3򚡎���S��e�q�nUz*~+x69��j���l����K_`M��>���:�_s	8a���j9�I}N�kյ #e���_S��%�zE�Sձ�'~�ҹ^� R�X�(����3W�+���NIG9[N�S^�׋�8�f���re��V�*�"��篜/�$�;+VC���صr]��(���zmQ	^+<�E���fE#�f]�}�;���Ξy8F:ZЭv%)`��� QDl=���Q+��S@\1�o�|r��jL�**���-q�Bb�.�l�'̺�M�� ��Z���^>Q�Z�7׿�vqXO�ܐ�o��=������B��)�E���.�u��2�� ���a�X�W�x5OR��!XƊ�?��t'�NG���qm�U=������w����f�6���B����]�	��G��^��ǂ�e��/��L���(�VgN���M�<�X��lh���%�����9�b�=ʵXoi4�:*^cM#�(.���Q+��43�] ���ޞ�!y��(G�?���c�r5��Fh	��wɌUkS���w+T	C�����;��^+�i�a/�Q��JD�S",��M�)���	:�,�����s�N�(�0���Dp�,�Q��4I?%Z�?Uy�$�ڐEU�~��1�L� �mڱ4�� ��wyM7p��!-�1Q�[Ո��"u�V�P*q��q*����1���$����#�����Yv�m�"i����_��d����'w����_����P��!Q��A����2£���:(e7�;�eN�h?؁��Ԉ%v��р�$�{5:�=@O�P��w2S�t�{�3-3B(�Bc���y���5�3��J*Ƌ�q3��@\�`�s.
x11�ջ8�ő�����]�D���'v��r'��d�z�5����U���B#�$kء~��(����_��a=���o
��<��
`byԍS�E�B�W��rK�M��
T�mz������$��j��\˷c\j���9Oޜ��E�#�!	^Z�0S��r�a��;{��ah�K�ߎf	�w]o���z���
��Ia�~HWf���	h�$o���P�/��ǟ��r��j�[��g6����08K�F�243���<O����x��jS�􁪶�-�.�>z7�.�й�Q�:���@zU�/�Q��8n엔��qf���
����%�uu~R�x��$���&��_�A�U��� �U���c�{�F�Y�,.��̐��܁S:���r�]*$ܥm�\Vk�"�+7�8k`�F4���a5����I|�F�x &�,ǥu�?�<��K��U"�����F��W�	R�#rs##|���'�\g�{!(�K��S���\��麟�����˟�L��w�)~eS�8?�D������AfU:..��7�5@��>���(!m�
�(C�A�/�2{��!�GE�E[ß�(DN7��z@[]�?��Ƚ�A6}f�oO~�����K���'V�e�pg O��2!Ϋ+�X���k# Vˮ� �=J�,���̵F��l�xQ�x�����}�"��z��&-ǧs=Fw�I�/�����/on=���<���q�Ku�R�R�JHN�
>%}B"g��]ߟg��˓(�����ʹ<�q�K`硝Ѫ��Q%p�dvӢ����N���W��	|O�1��G�Q	�=�,{�M�/Ķ�"x@�qS�����x�T��+����ѓӪe-4,�y��c�.�6:Y�sMB$\�Z]���J���/0�B�3WbJ=h�:	�u�tn���[c�R?�aO�� 1�E�Wra����N{ӥR�
��UB�K�#|�3E2��TS:�0%wQGW-O�+Y�z�n}�1w����+�@���?�䖹��'�[P�[v������x���I5v*E���P2���nmL��ཡ���̀�`l'?*GG���(
=�F�9�}pF!�4�a�Ak\�\�G���{�Z�l��ع��9�lԫ����LR���".��su~��º�v&Ԃ���3Q�Ni����kƾD�YJ}&��t�S~�'�܆w�l{ƍh��1�qU7
�?S�+��ti�9ϲ�vx�N
>@2Vn�Z���s���t��:bz��7�-&\�ɢꬺ�����!	�@:=?h#N�wq�����6Wy�X	�|���;s���NIP�:���<�+�&���b.��m2'��݆��,`Q�*��N���;��	+�����`��^w���5J��9��xտ���ܚ�,K��]���hu�<a �8R'���x����y̶����?p��M�i;1��$v	���9�,�آ�%B���2�R[.�OH�_���u0����ھ��܎��:ίO6i�EI��쀚�b��1�F����D����	�˥���?�ܲW�Um~k���FϩD��'��9~|c�`��13T݁����Rz?�K�MWr���6��H���E��^b�x��U.8o�i���D���ϭi��Y��,�����{η�&��n�j^�*�7�pZ�z�`���5G�;7<��X�Ago�*�aؖ�����!r2��C�Tݫ6��%%i�$Tپϥ�iu"4�m���6܁�X�b�����O�j~�����bdMw��a���������G6�����⛾�>aET[�G$�on�8X�_�(��5}	�U��y%����V�s&#2{
f��ﾙ�,�Ҵ9S������ĥ�9:�V�ܻ�\�+0�fx���1F�=C(��4�x%="��x/��݂�5΢�Z���ќ�4�j���>�?E��W=
M){Ard��!&6��B�W΄VV`�NT�(�:5�����+>��잘�a��븋�Z��l0g�Ơc5����S�hl2V׭g�ݮ��x��+2�x�Z�#��j0�V�9ش�������o}�W�~�|�?Xl��z|�B*٪�oR��o (.*�Eͪ�띮�}����X�`Z�r��b/�3a9u���޸��#%D���b+;s��%T��~�W�d���4(�}���o5X���W��-���$[X�V�W.ے٩r_w�r�\�3���dPU��V��$��L#���,H��i�4b�F?c����b�������z���q|d-#�(�
Z<�o��p��X��o���l*Ԥ�@���P|���w���,���S£u�����HX�P,��Z�G<�1bŶ�^�{f?�������a�����dt;��}^���$g��Đ�|�hX����"S��w-��;q<V������ɥzp&M~h��q̷jsIv1�-W�m�q�87%X�uht*���11���(�k�Sq����`!z���$4��8�e^�%�����0���*�قv�Rwǽ��땠��v`�ٶ�cg��C��'�/�l�¢j��&��ǻ�����_o�h���͠�VV�%��ωn��Fz�P���b���L�eB+�$/`- �,��;�<_�5֡? k�^�{�m���O�Q�]d����^Q���;)obΫ�S�9#<�c�H��e�F�_J���h��ȓ��;�ߣ'���F:r
3Ե��}(�c�|�=��y����+�Ho�[�֑��(Õ�&dn��&-n�&d����\ܞ^� �[-*�d��TS�+o����#�e|>����)������t�M�y�f�t������x�ۋ�`��K�д)r�+B��e��lcF�:�.1Zzk���	��ɏt�a�nTC�J ��~�T�ި��GT�mS� Q+���*UɆ� d+h`�MɂQbtpؼ}}ڥ-e����P�-k�	�[eejhi-I�1�OƬ������Vh��;6qx�[����̠ၶ�E*��1����-P�,켅��r�T,^�U2B�j6s���AٷW{�k�+H�s��l�h��ڕF�M1���bK%�F�(1�b�e�(��䃈܊2e�#|T�UG�6��F��D����!D�?s�t0eq��2#k�2�k	F�SuLc`�U�!r��ֿ�4�;�wF@lN+�H+ѧ"m��z�`=�*}�6*�O������Op�Z�E�+�;u�4B��f��>��4�!5��
�
�^��$d"C����?�?�_♝�W�u�p�	�p����7��T!4�v"VK��Z./
�/��j\�;0��~Z3*��@��a7��[r0�`r	�
�:�����z�AUN+�s.3�R��.�^p��r��}:�?�V�
���B�<ܱ��)�$UXۜx�aU&����2�{Y�ZI����r��x����y���h��Bk�?➯\׃i܎ߓ��nHKDS�v��8�h|��vp��&�>Ɨ�2wu�A+?'��E1x��r��p��	I7��=��G�to��(�d�6Gh@h��g�O�PuVk�E�|� h�{�34�#U�g���*l�:��@%NYpTc=�N8Wc���ˤ���,T��pF��6$	���7ݐ�R��2*j�y�2�(��cR��(�$���0)@�������:�|���pn�����Q��"~���ʉ$FM巃��1��*6�a�����c�`��uMG��^�i�����*����:�w���>��5#Ԙ=�cg�Ppu|ף�s�H]�]�aO�d�'CR%�p�EYf�!Dr%� t�C�'�􉿅D�(cb�̐ x�nY1O7�u��קB��l�Ƀh���Y�3/-
p8�ս�����(ը�������"@�L1�6߯A�*�O��rg���� ��p����z͡��ņr���Kٕ_\�Ϩ?<1��_�����<ы���%PR.�B��ݘ��o>% ��'�����)V�`��@��P�)W����\|��J�����d5�z����$�g�h%����T����9A���C����\�{[S��{
�q
r6ĵk�c�������r�����C�ˀ~�ZAJ\�1@��Ȝ� ($�p��P�
� q!�FD�z�r0���'���H��>m�����f�џ��^�G��=)�%�kf�2�a���º�l����iG���k�!q]�,Ѓ4 ������$�G��d�Q�:ZD�V�4/�	e�>I�'S�r�rA�aԦ��QC��e�V�2W���]A]`��>�PNIV�k�^m!�.!��Zf�)�Z��=�^�<Z7@�#�& �a���� �[<@L�3ӵpPb&[���c* ��55�[{�]Q ������S�L�w� Z��mi���7"b"��4Dˡ�eѡ(�NG��L�M+{���T�y���G�A����)������n�\b/;Od5�"���z��>�8�{�Q���A���W���!�W�w�;�=�& 2:ܚh\�l�@��(kt�E��Vh�.�.4H�u��"�|��}ܬ��:�h���)Kd��<*P%v��j�淩�4��l�!dg`��]�b:�����y��7��"�n%[�m�h˼�����{�Xc��J� 
�d���20ѡ��$;%�PpAJ(���
*����s��r��8ni�B��X�cU�<�ꫭ!���K��vt+&�:�nl�Q�٭�?t��*�pF�����{��g��~�Υ�Dgq�a�X�n��
�N�aL��/�C5�z�l��/=K{\oD�cg�v������m�ګ|�v(g�	Nwf�� �D/��
8�M}�������P�iT���h.�~G�ѱ"ˇ8.Gʅ��n�~j.&S�p++�K�x4�Cb�A�@F���j�P�^���/�R����5�gkE	{���.K2��?]#7���51[&��r�bԥ.���:��i�q:���X"*�& �TǊ�L��T�ű.q��s����a�@��0��w��(�X�S�{:J�'��|�����=x)�l����%�����p�)4�α��2�;׷�@3��Q4�j����Fݸ=�R�S�BRd]�#��u���� �ɫ��a9��_�?��$�H�`dk4Q�l!�޵N�`u������f-���Э|v0ѭ��C��tn)�1ڻ����i��(��z��ش���;����5��H�dZ-��˂O(����(�h���ɸHG�R^�����o�?cMj�:M���l��1lI5���P#�Y�|�"��k�>����?TL(�C[�!�`�Im	0Q$`R)���ɥ
�F�4��Q�����i����:$M�;~K	с��T��%v�ٵ��T_�<�'T����Ͱ�dlp�O�e���R��TtP��O���IP(��
�a��1�!�Mρ��1*?�ͬZ�%W�AYO�v���f/ͦ����T,3@�˷��&r~t.t��C,Y�:�U��,���F�:%���mR�q��T;��@.4����xRtu�d�4���W����Z�|'��F�k>��*<Xn�ƍ3Z��O�3 �Nn�)�Ly�u�t���,s,s��VƩp�Z��R�.ꍹ�����s)xy�F�̋s�濥n_
|������hR�)�i�J��-��;�꣋�.N,1X�W(>w�9osW�SxU �V��?q&>ț�����h��LnO��E�, ��`Z�;� �h%Xtp (��V��B��i�cU�GU�d�����o�
�
��Uf��8~�6f����2�i<��x.�b*��!H _7�ԃp8�A���Oi��6��l�E�j�K�3Ϟ�ivy���^>�f39�Q���^Om2�	Hp�j�߱�U��Ο%�J?�ƯJ��)����E�rʶ� �T1USj��d��H��̰L�ۡ3nO��h���9��N}�� Gjqϟ���idX�Q��2�UsZʿ��f�4�� -s��=�zko�=l�<���x�@�oxC�\-�E���l�da������/���Ry"T���a��*�i�90Q���.���d�%�؈�c���|��u����=!uKL�$�����V
�����������|i��YNP0�������cT�^+
:�Ӕ+ M�
 �鉋{�m���$�n�C�	���j ~������T����XN�ԧ�O;F��'��Ĝɣ�ߚ*�d^�Car����r�;��R���A� �  �<�+]]�2H� p�Y]��������+�8`����C��������Aӎy{vJ�qn�2�\�|
w+���{������V����^ LY!�O%<^O��I^4����W�?^��ߍ��ܝ\����{31(��N�7hmrQ����:�.�ԫ�'镼r������:�n��J=�ĳt��t��^�*0�dV-�'.�p����֛�y����S�G��Ψ����͞����hEgcsu:��+�@t~�Fܭ���P%ÍQV�V�l� ��I�np�x�s�v��q�PW��ó��T8��%!ɛB\�'�qF�tz<�xUq�"��Î�0JQ3O�[0_߄�|1�h��D�Y�
�
 ��%
�����9{~�k���Q�8¦����F!c+���K&�[�²��,�ąa�ҽ`9�B����Ö����$Ÿ�}��X�E$g����_�#�'x�whxs�R*�HG 	��c���#M��Ky�LL�ͻ،yU\��nB�Mg����kn�b��%�f�x���So���?��nd�>.]o-6�[��������<�i�F$z�ӧ0q�L��1#�D�xދp�,@5Ҋ�ڜН+�=h���'$�x���\BR�m`Gb{]M�8>��8K�j ���C�4߭��Ε���A�y���/�n�b��BҜ1�U�0l�����H�Um���ںMI�.�$��S)�@w�8�A�W��j���������:�y��
�*��hWD����b�M	S�^*c� LL�ڲ��)\CG�h� 
�؈�C�f~���|��'�-�k������ޕ�j��'
�U܊��-;��A�]����k��]BZ��.�qp��z��RM"
ٖbd�S��I�A��%�-�eG�L�ț�H���`���J�B���s��܈��J%(ToلN^ �����������r�h4Z��ҝ �Ş��2ae5�+�;N�}3�nv3k=��2]�ey��+�DLc4�+J��{=��,#_�JYEefBJk�(�[�oI�Ζ��[4��}��>�?f-,�h�	&��%M͐�.��8U|.1IEv�"����{�:�{_��6�o��Υ�����'6�=z���tI�0��G@�yl�|(���p̗Lo4RxEE������`�M��|��"���3%V�=Y��O0�-P:�������-�Y���a��q��+~���ruśB���e��ǉU���2,��]����'O�����\�P\�Z�S�Q�G{e����ޓ��7��|zh�4 �tѕ�����n�:����G���	27)l��T�N�[9ƫ���%W����y)*p�ݷ:ʣw�%��_��&����G��\�Z9�qq��r��c�~ZJۼ���z,�5 �s�$hBQ��T���"E�O�Q��qfa�`t��BO�Y>@��ٺLN��0߽6��a|�ľE2+X4���#�;�xT�y):!=	���N��}�=3mo�c���@�ʗ��p}wy^f��,�P��<M����\5�[�o�������-��X3l�~D��GiM��O�i� �=��Nq�	�y�8���|Y֎K�ԇ�9Ó<vW�_�_��le���s�]fN�
k%��%9����)�Uy�谈�2eo��K�_;�	5��1|�)ΐ,�~����g�����	�@nM:�P���|_ƄI<S��:t����� �LQ�[�r�����(�A$a������2�d�a���
����s�����F�hH�Ոu5��%1j���I�[��gX�He����g�ڻ��Y�V[a��ZS�9jPg����)��-�r҆���c���ĭ(>c�oL���Qk���x�4^npק/A��e�6��,X&U-¼_&S�r�������8ؓHk��/1_j����%K���+(Dh��b|�C��A��G�m����Q?��7�/le(Δ�]𪷓~ܛr��UZ2�(Z�hW�q2��Y03���a.�K[���%��ڗt5���Z�z��@���g�9]K]��.)�����b�eSU?�J���t��.vSDa��^T���C�ϰ�\
'я��WAq�&f��VJ!��]�T9tBf	���S�Jg^G?� ��g;����=�.[�3 ���B��=�w�Tu�/m0>㤿z�1�\�%ح���޵�v>5�=f���	�d�L�4Qb�U��*jw�-��0�����#"�{6&�w.�� �#Xm�����p�O��0�#���g�N�"j�+c�^��m.[��BQ~�p����������j�ϱTlV1*8�D�ZJ�,<m���Kӎ��`�,
؋t;�� ��"���@rK�7���
��+)���G�����T��Q�jmKh쓧Sӻ�&�-}|f���-��B���xN������>�`:��5���mf�Q&gJ�0���o�wc���ϧ����̄���**_��E�XJ\jX�'v{��r��ng�b���(��n���=Mt���	���vzu�՞�_�*�ί�O;k��Օ9C�O.N@UN��E��rD�[���~��J`Q�Un�$�f��m7l�6~'E�;8f�]� �C�O�֎��X��M�s+�!?���(*Æ'^q���"nb�b���� -D벎K��fj���U܅�b����7���Go!qΉ�*
�Y����k:�d7�0i�����ꌛV�2��~3�m�n-t��#��PA���Q$ #l��8�Ѯ�۾�B*%��D2���І�C/�J��f���f٥�]�V�c��LN`�9t�!��H$yo�*w��3��3�،��2H��h��'���;%�`n�֣�=`�D�)����ϥs�	~7�^���75-��?�y| Sp.�j��X�Ѽ��	qU�Q��A��l�4+��T�용�P+*/���XB]�8\�ZK�8��]��)�7�c�;I?7����-�e/is^���܌q�N|x������*�Z��隡�����q��%
T�2Ծ���ت2��������}��D��Fo�U`�0��j�X7�Lk5�B�¶X'�2j�ɘ������@�fA:q|�u����z���d���T�v�9���̽�d�;������c��p
���v_�ư�Iθ˙Cx��-;��Жl�x��B�#�;��C�$h�Ț��^�Nξ91JZ�g\IR��<K\	��kM�\��F���s˦ pG�~���Pt�T����q��?��Y¼mr&f�vc뽞�-�ڧPt0i�3i|����H�R�ྌ�Ħ�5$�<25o�(i�&�򴈧	��}���.�[�_�V
��������#�[����o����ax�p�n��`:HQ�R���+G3�r�S�1iab�d?oqj5���ßQ�x!Y���r�T�uծ����6���W�=�'�Ԕu��p~L�ތ$~�ɇ|4RE���:�0�#t��"�xy���#@��7[O�]Q��L<�]��v�2?O/��<!�MX�1i�O��=l�ޞ(8R3J��D� �b=�B\�#Ie���,���<5�cI	�\�I�,�����G�?r�����IƐ�ϓF 2;B-�uć�b�J�}ħ�E�6o|X����Ghy�_1�H�ČsjCI�:i�Os�k�����7�3���>� �����^^1�+����%���Te�V�N_vw�}:Ap��޳�V���WF?Q�#��=j��+:�Jy�̭�b+9q����&jO��jl��1%Zq�ٍP��DK��D�DG�c���1�P?�D`��H!ݞ���[�'l*ʷ���{R���-��ԓT����tK�&8��$��k(�7��nҜ���{����o�a�N�uճպ�Lg[�w
��X�}����T�k�4H�K�d������µP�D� l� bv-�5����~�^X��Д l��ە��/���
�&��ˏX��:�Q���č_+u�z��o?�����\O���m,��UE#�3)�_&��,񣒵���i�2o�kؙ'*�o!@�k�BJy��!����.mOA��72�c�(A�p�\��_iNr�A��B�l{���jf�涤'y	+��R:�='W�GlC�w���%���>�X��i�q紮���J����]��\�Խ�b���@5Sz#̴9'A(�%!aA͈�F��؝�dk��I�������Ӓ��m�3��)ܱ���?Yy��?�Y^��R
U�����Ȑ��81��I#|�c�V�3�Rs�h��#	)g�e����s �g�����F�
$�3p7!�#��VB}�q�3�6���[�)i�'�y�q�M���N~R�Xb�~�����{��Mo~̵���gT7�q��f/��.�h�2���8��"*���[u6�B�b�x��w��.3�=�!U���>M��h܈g!���@�<_��E�n��c2���I��X��}��Q~�H��w�ȵ>p͢���s��Q��v���?
?n����Sb�q@ax��VS��і,q'��p�����/	0��N |!G�v���J1�ٟt+�-~߭X�Q!�W��wB:�9c3�����'��?P�:��gT"���Ve�	%�[�0��X.T�e��\j���!@=��M_C�����nd��Ng�������5��q{�²auWW�߭�q���>����ԫo�L1���z��B��m�MI�<�z(Q�@��<�j��=�w�D�|>�]9��e�{;�n�3:߾`��%����>�C�^�����R���Ӟ�%���6��n"K�q��'r���x��.E��\j���U�)"_�p+���W +�r�{bA�G�i��o�ۥ��ii5+j��+���#\��J�
�TH�N�CiAx?�`����5�4GI�o���§��s
e�SH�LNP���y���!C�O������CywNv����\��翗��h�)ĞZe���\C7��P:�7��e�RK�⚏ϒC(��/p+uAYV�fB��of��k����Q.sv�
�@�*��^��h��P�� �\�5Z.^1S�AK.o�\\(E�S�~.�^�M�Z����H�4#�kL�E�Ď�Q:�90��Z��i�㖣�*��o�hp����	�
QOaWu�h�ˀ�ׄ��}�e�T�3�Q(&N �^�-uF�n��)ԡ77>R���au@X��R�K>�w0������|�}��Bw�*�q��3)��
���<Ǻnm�I� ����>�1��4x�����x�����փ`�t�V�H���=�����{����i��U��r�e��=AǺtc�4�T���O�ߡᙰ���� 6�(�5 �"Ξ~ЎE|n��̹f3Tܳ��ރi����H��`�S�V�+g�a��A��ƹT���I*�3���{�����`An���)��W)�c,�xC,���ͼ��cL�9�I�q���94
��%@ձ��@3�gJCC�B��I�{��u�ӗ�B��i,4.ܘ�륗QGf/�9ٕN)��9R���QD��؇A��գ�A�E^�ػ��8��+]��`���/�*��N3��ъ�]���`��;8Q)�Af�/��d*G>�R��H�hGEeoq�z��8���rC/+�C�&�������D�)�q�|*�~��k@��>i�X�b��l���vD������v`�~��R$Y#Q�����4\��(��4�"ע���[�����jW ټRU��b����Xfb?>�������꼍�c%�C'�;����+1Flxq8�&�X��z�L���G�p%�X|��#TSL��|��LL��	�^�5��r{�Q%X�MF)��q����{�Mݺ~�m��D?#��8&�r�/��FU�� U�U�)�������"ޞ��^kS�ش΍̲H������d=�t�#q���9���6�e�=3��¯��N}��5A7j��������N�wW�l 6g���u1��Wo�ڽO���CIK]ҍ4HȀ� C	ҝC	H7H���
CI7�!�����|ߵ^��?��>�������3�Ԕ�'L	)$L)$��uD���2i�};H.��h�{�-¡qזE��9І}s���H������I�E���F�����ل����Z�݋$��U(F��'u'�F�G^��������F(fHY#t��Ϝ�KM��K�b>��Ѿ~��"҂�Q���.1�L|�s����%��?�oUhŷ��a�u�މ�@/8E� `��\W�j|�gz ��;��²��0Ӎ&��#
�09h�ûTlAZ��ƞ��՚��;���Zws�>kӧX���?
�L�c��������#m~S�����7?�K!iERĚB!�V`�G:L�;ߨ�YX�N�����@� ��ݯ��jZ7O4:C����}ͭ�޻�왼T�g�J��E)�@�/p9��v�8����#y��� �c��v��U�l�ie�P)'La3OX���.tR��!7q�_�!��T}���vj�`%�[�y%��o�i�GZ���;�ՋA{��s�
B{z�_B�؎>�x�CEo����������0�����C��-΍�/�`dH�:R��'���06�
�ӿ���n��f���Ă�������7x���o���*p������t&b���-��#���щW/��OeTwy��rbF�1���:�@e��~Ar��q�󄡝�h�x�z@��\�'W�os��3ɰ��Z����^���Vboq���ǅ%�d�"O�>U��Q��#�4�%҇9^}�Yu��;��ld.E;��p\h�b��g�rbm�r���=�z�r��W���{�Z3a{Y��Y�B�t��P�H/���\;��9W�H�o�������t�� ���g��][���0��Ȳ���8��m<�� �=?ܤ��
�c��;�Cv�T�T�����_��=�-K~�,ugP��L�k3!]S�!�ޥjK��WH޺X��*5�J~v£�¿*@��+��Kһ�B��}�t�` �Dh4V�/�����{,�1GE`������"�IL�e��vPB� *��}阣��<�	.�?>բ�B�H�b�$Z$����J�Q�GX�*i i�;3�)M���K(�.d^��\�5WV&{��e��W��E��L}Et8z3��PX���;�<b�;���	�i�԰L��gPc3�G�Lt�{t������q�Z��B�/��Mw=v��9P������xP�[�x�)W�#i�j��LK�nU�]�ݦ�a�# sD�Q����w��e\刈?��vd�Ji4���y�E���NM�뛱�M��88n�dGLSY�7��7���j&��j�Q��/je'�Pq@Bu"h)�Cyy�����*�ي1�w���
�w�bhQ������g�Z�`I��O�?M�0f&S��Vxo��LX8���>����;*Z��7���
���,w��n����W�;�9
��/�>f�@����O7����ɿ�����m��ラ��.��Ł廎/M>�nf>��S�o�/ws�a͆�d<yl��P��:B��7~�U����5�
�*�Ѯ4<^Ut�e�4[�"1>�.��eq��~B��QM�����ԻƩ�w̹QP�j�U7#�X�:��5J����ނ�Uś�H��-Ax@�6��Y�)�,�!r4� x�y{٥dd6Ar;��)�z:����Ib-`�"��S�a{W�����̀:�Ռu$aa�Rq�0zX��7�K8�� �nȁ#��m��GY��{��N�]|�G*��\XZz�ʞ ��G9YeTѣE��(���g~Dӣs�9tR�
��uR�~�?��9:��vYb��2�������FU���K���ֺ�x�
DK)=ZI��.=}�����~�Ҵ	^H�X��`��9�3�-1���༭�1�X�Y<�y9L]x9n�
+��z�ˏ+���튛g��
�N'�3���x�cV7�dg����xv���j��gd>9FIT�L��ൻJi���P���!���ۖ����'��_Y�����I�^�s��H	��]&M8)3� 0��u��6���$Jl��bf
��_
�@��ˍ`G<�۹ń.|��]�����5紕�@���J)�6j"+j0�:! @W�F��|eh-��G[�܁e�rv�PT#�?	oP��uɔ����r8V���T-�f �b�$��E)���5\8>���ַh[�ff,�N��we�9�p#�qА�����|�C�C�*Φ��H��|�>�#�G�f�k+ ηt�i�q��E7|N0{\��[A��.���	�XL?�[ķ�v���W� �2�������˃l z �m���l�	���_�$9�M'��HC�EXRU�����~=#OA��)Q=CϱD�AT�GA�/�u�o�OH4�*�� ��LGJ�n@��	r��7^Z�pY"��2t3.�	Y�Y�GQ�����Cu���)�XjHhvky�,S�rr�̀�+�S+��?���5�}����v	�&��#�s�8J����=p�4�� Y��X���n ��:2����� �:���ӥ+'G�<+V/S5!q	�ؤ��a:s� ��|��p�0g���� =k_�#qF?3��DJ*W�z,��r�k����!� D��#b����qq_bWH�uװ��p"ї���M��L@$��tDa��!Y�A_�r]��3}XW��mXjB�;�
�U�;�ߠ��O�Tt���d<5b"��DQWStr��\$7~k��',���pU��)�X ��.� 3!���d�������H�na���F�
���� AP�z�#NF���h1/Z�j��:�A��w�u!�������1xm�ޙz���#3)�?[������/��@W �Ik;4�E������
�sU�v����U�e>D��n��2'����"~��H'�_�e���3�)��>c �<���Ǽ�c��AE��+�$���c֤pP�]x��]���u��%�b�����dj�m�}\����0��08�����_"[Ym��T)����[s��B�o�q��A�I���L��h�>:���LR�̈́֒C VS34fT���J�v����g�bix���F%���A~V}��"n].-�ޕ3��~.Zp]�R
R D(b���~�jJ1s;��"��*#��Ik�숎���JW�N[0��߽{�Qj;��j�ZLi��rKy����zс���G�L tޟDp��x\l�/�Q$x;��׻�-�p2��{��6�0�խ?;�#!���g�1EX�a-�y��`:o�P���6��"<.��ޛ(z�w��eZ6��C@V%��ۍO�gO"8Q��Ln� v����-�������+!���-R1C���>^FQ	�t,]Rٌ�l����NW���T�]$_�������<��ӊT�Tj�	��L����Ua���p�ꀩx6�-��:3'���WŪ�1������8}@�6�籜�j?9
�w���o�]���ś�eSF�qI�0��]���ľ!c�i�sE�ԟ�ʊ�g郬f5Z��v8]�!���c�k㏇)��u3��mU"b������ �t�<=Q�ʈa}�:W,�N#�
Ç�srh�������BqI��������}.���g/�1
�fׄ�up��c��]'n�AN�/��72�EZP�a�����-�-�� ޷F�=�*��f���[�4��g�.��:��.���N��E�3K�yx��Y�Q�7�FN[�َiϣ�$a�Pj[��
��9� i� �=M���:E��X�K�Ǭ��]�<��zj�Y�(jW��������J� �vq��Μ���1YW���V7���ه�ynR�зB
"���J� �Z�Kp�0~-�u�.��ʏ���Kѵ�A{�����$>T?�U�"��,�%)-�6���ғ0$!.;���D�j�bl�2��?�pA�@}����˂�_��#�0����_����L�?9�ʝ���|�_GZ����j�Η{҇��0`��N��S�r3sldG����e ��w`�&B��F��=�\Mg0��d������[�+R���� �P��)�'�	��!�S�����+O���:ztY��;x�K�ޭ"���͍kB�CK���I�f��9�RBem*�3�Ӹm���wW��s��H!�U�G[N��3��# ��`�r&�o����/�cl{�$�����=�K;�y����/E���
��tC/J޲.<!�ο")�ep\�~�$�	�~n}��ďL�XI��C�:!� �%r��:n�%1��|�8�^Cђi@%��ˤ�:�;�3~�3*��������|��߉������*Q��T�1��Ź�r�� ����v�L��(���P��3M	���S8�^$��|,Z�+�g�X��P\l����0;a�z�i�g����"*�m�o�a�oJQ�d���Ȯ����������Ӛ�U���N&�;�j��}Ō�[|��/J=���M� ��L�~���U"ѽ�JR��PiQ�'0��N`�Ԕr�^"
�b2vՖ�D/�)��X_A[EQ�YP��7=��\1笆��$�<�H�`��7�bD��xӣ�7�����ba @l��
B�'��+T�Tʈ���Q}�H�ܿT�q�=���ba}���94'#B�{�#�+�)��M'h����䠷�a��^��=���)��m�QL�A�v�Z��!OJ��%�PU>U������T�nQL���^��,`�Fց��>�\�Q��y�B�/<��1X���]�Y��C�st*}9��ڧk����ߐ��w=Mbv�g/C�}Mǻ_;�6�cm̬�W;��:,?�4��Z	$�KV�����_��p�~�-#o ����=i:�mT4{�s����t_�g3���J����=��D���t�1�'��@j����o�d�qS��%�H.[�F��:b���z4�1������`��K˙��OL��"��T� ��ͥ���2
(/�a�{ݞ��&x)��^�1 >\�I�����w������~�� a�0|H�)�Y|@D���m�w�r���t��a9�>�@<z�������!�h���Q�J���tl�*�z�I��E(��j0	�
��` 1}3������o^5��x~e
͝n�v�6��7�x���GB�T�}'_��Xo�}�t2�<q����i��'�I�`��Rၳfj�@��*�I)+�&�1����=�_�M�m�T��d&H�*���)^��e�8{jP��џ���I!��N���srt
ݳb��~Z�$��?TnU�
�NƔI$G߮~3v��Nmt��γ�Mb��T��}\
��0IđO�]�|�W����e5�
9�l��3���e��~l�)3�1\��q��ƹ;}&��� P�f�� ��jxۙ�bV�D�s�:2�k�g]�ų-F��ު@�kה�|��p�Mk8my���b���qm�$����ggS�M���_��\ԅZ"n��3#��9���)r��H���/b��
p �^�=�D�N+�X0~A��5��T�NnV�}$]��Dq�G.̉G.�JF&����-[�e+[��|磖KY����Ӊ����G��o
t�|t7Qr�q^~�u�[[�*�!��o=�ߙ��W��d��^[�%�����a~A���uS�V�	6Fy��Q�i/�T&���!q>�8,[*hE�/q]
��&+uFx��>�qv���4┧^#�w?+l�$���e�4.�.}�aTnG����Y�R!���<�-�
J4��{>J����P��;��@�Q�)�]@�� ��/9�ҢNh'�I��i2���t����N�p$�У�Q��8V1�Vp��e�N�~�J�~`�?�L��e ��)�+M �^� �g�/�y�:�3E~�N�)"e��V0ė�[���I�\�.D<�?\�����>�������۹s�0ѯ�7��Lg���b{�������	��_-/���R��>}��W�#�u�g�H�l�&�`:�}��|׶��ɍ?h�n���0R�9n��d�1�z�����%�P=>f.!���N�<�Fy;�	~�R;�����nx9�n�̷mGo):2�*�
T��N�x��Z��ϯo~РU	XE��ys�yzydN��U7�I�wT��3�ʑ��U8 �4�����Va�t0,��E5ՆfL�LH�I	݃S@5��:�ɦ�*LM����;J�w����n�p_H�$�&��R`�b?�����8��R�{j5�T���a��/l,b�� 2���Eџ���j\tEo�����_/��(�����KJ9obC���5��Gi�fd��59�>O��/�L��2o**׈�L�+�����<V�czRs��^gH���,a7E����n��Ӡf5)�`��4�����.<�sf��Ę��(v��6z��F���_����;�+G)ݗ@�R����L�ˇu�/h�把T��j �e�w���Jo1�c,�'&}i�7{닏 RYW�A�1�zGN��]V ��piٔ�▴]�����1���r(~ݟ@G���?W^���"�����	�M���A.�䙸 ��	�8�o�Y��o�4ӊՃ�>"S' \���ͭ�!@�!��C�6�-o�_.��v�5m����<mb2�Z����8����K�2;.%Θ�:1s_IM49�k����z��]�4R&�����NA���>�DF�s��Y�( 6b_� ~\ϼ�=�X�©�}a0q��R�S���e���Z\80(��çFo�q���Ʃ�/A}��:^t�����B.�Z����� �f�s�@Z*\p���m*�v�����g?�1
�T�;%���2?2TL�G�H-����윲�KÃĂ�TzK#����K�؅���CWp.�F����:3tg��'b"E.���	Im��ؿ��7=�i����-sk��u>�P>!ksO��^�����2D��|@B�<L��v�{��[�5���'�ִ�*��=�������r>k��Jp.:�}��휦I��%�ڗ`N&���͕��ez�YB����	2���������X��*�vA���y�����5~.��އm$�U���
��HYʱ��R ?/w��L�����]�&vT�����X9�ֽKL�/�]$�gn� z*H��4��-���?L'�K���P��^�'\�?�>����	R>�|.<wE�I��C@T�4�(CQ�Fᴤj�����XFС{$)�r��o��R,�&���� R�M��(n��ϔ�f��txQ�D�Pz�G� �G���b%�ٿN+l`�)�Wwل��6��8�C�[(�B�j��}�3���l�F���!O��Xޡ(���kb��V+ҏc�ЋI�7Z�}��B�&��n��R���ݐ�5�k����MSM�29e�4�͓m�E�E��/��w�	�^حUi���Üi��i�d���
�p���j��l�)�MȾ��a�B�u5�A�����s����i�z������ڝe����8n�3������@ɟ�>��F���ZuE[{��M�n��w���E��G���Y�|>���ґ��QN4��'��4��gR��q�3�PJD��K��BG1м���9��C��/�ʭ5��G˘����#���$�KA3DP]?�����
X+�f��'
P-�>)��Y��(�D�Y�^�a���r�@�3�KҶ�A�hW�j�)c��a�5�u�<}��lx
���ViP(�y��wx��_?j�P�9l� ����?�k��7+Ӎ���3c�+Dj;�-��'[����c׽��Z�Gj��l]���X4�����GE�Sh�E���?G�]qs�2R:���� Ռ�x�'��X��k,E� ��ih�֟�9Ӷ5��&pqN��O8ޞ��UhU�0���s�=xiE��pM�����n[����F���.!���M� ����s=�'tt�2,ir���ؿ$U�X�N�~�������C`�,��>&��z��4�'�
i.�K4{�ha����)'&CJ�8	�N\Gq��Sh0Ć���>q�������ߺCs��E��
����Y[�]�BQ�K_��5&2T�d	V�#�$�b���w�ϯ���ᰶ�N��K����r�Ҟ����"�5,�/6A>�>�o,Y߸QR��D�~iQ�(
e"�k̈́�z��
5�L�1�P��c۫b�2��f��y`��=b��^��^T���&&�,�_�:��� `#p�#Kd�����ϸ#]Y��١Gk�|:>3s���4v���P� "2��w�I�ӯa���u?
��\�y~cy���J�@�V~l�Xt�E��G'X����+]� b|,f�����V��9%:'� كq`�Y�qA
�9�>� �#x���C��M5���a��	8���<|��S%���)Ǝ9AA���nH� ��o
w�����)��m���,�S����Rw]��$����~Kv�qk;ߑ�m�8�֓�;��$q�����V5,e�n��H*��VSF@/��Q��*CE�����/�s��P��ź�c��l`���d~b�O��Xl%�����Ŕ���V�����5��v���T��gKD��#�۠�?ե�V�='�7 ����@��ԑI:��Q���m�So�L������!G2M��ݿ�P����sq�����f�2�]fO�ғ���<As��\�����sv����h��jT��*+��F�A��P;�[���=�P����;![eG�1Jm*0E�P���Y|G2i� \����ַK�6�5�փ�Xlk'��?�o�+���jj"3�3Z������a��(sG���79��A��rzY� :�T�Q2ϫט`(
���?
;�>ջ�>��k=8�b�<��*9Y��{�_e���X��TG�N��NW�4E��aS۠E���G��V�6U\�Ys+�� �I�s����?����V>�2�D�>L������<)[$S|z�,����g�_�d�1������*�~����zD.�~.�h���X���UJ�d�USi�u�P�d�P�I�4S�~��R�ѰV����խ��ȭ��PG$nD�'�b�i*:NU�(^��)k�L�b۳�����)�xT������L)ɠG�è�_�J&������z��i��\QErn	���h�4͝���C�4�	�V�f5R���J@B��-�����C�&��?�<�Ш���* �g�]���["���=���&��?a����h�F���vǭ�L�\y�F��ΑC�Nq���� �����E�Q�C�"�)y�qS�R���h6�Q�	?�XJ�v�t��7!�n�1�MN��_C._��lnN�9W'���G�ۍ������Ɛ^#�B�
!N�ܟ�+*�T��W���[�*���+G���W��5:g�˅��]�������~U[$p�+�)�l�V���.�y�++l9�&C��Ľ{m�c����|�xŸ{�
e&�F�U��#���DW-��i�9��������u���?X!hƋ=F~A�G���-�bl�>9\Z
b���@��#���Z�ll�]�1f�����{�|����~u�w��������&jK��Qy���d��2���˃�������ꖿj9GG��<���Y�����[���Zq��A���FCՉ�JK�;9�O׎ּ�OEã	;{�m�W���~��	ͣ�<�$R�)�^��4*��?;m��i{>�$�5�6�18T�Lq�V�@KO�{��;GҫR��G���7�	������{F� ��>�vs/���Rσ ���dve�΢�tL������� Tj���J�̷��]O�D�¥�X:�3�G��~�`�4�В���B�A�[�����&���kI�b�cu��I��)�|����M�^��
�/�,��ܻ$*Z@���g���:����I߲�8�孭_
~m����O生m��>����_���o��ء_�Y�*
�Yer��h8���q�c{�����]RF��·���tO�x��7v塑/ȿ6���x���O-�p�T�YT󄯊��Ô����lu�{��M���ʙǩχy5��>4x����I3��'��(T�h%mI-�����a�Se�j`�@zcXb)��4C�Vb�Z�.~���)�Y���ն+ҫ'�=���� ����� �_�O/�ׅ�bX����KZ�3mm&�Ֆ�Ei�mH�]�	O�)��`��������5��;9�D�ݣP�$�ovin�u*j��=eB9�)?�tK��Z�P�b@f�e��ߓm�k} g~��/�+wu<yt�=:꧝��V^��{���l�Z��ȶ���Of�os���h5T$�T�@�*)_r4/�2��G����d��z_���f?7�Qz)������H���P�6�l�J~�|�g����-Y5�)�ܰ6*����f������ ���]�1Ϝ8S%�J�g�x�;Z�_#>��sC�ZK��s���i�C[�ţ�u(Z	�˚i ���')fU�9��B =�ƂiY.z$S�G�<�F�Nrx
��E9 ���r.�a>!\Υ'U����}-b)Χ(z��<��|���.��X��V�L��JŁX���o%b[��k�/GI-�f�ũ2<v*Y����z.��v6�+�U|��w�]����6:�͡ܦ�}F�$rg�L�_��P��a�H	H��� �GZ+K;M��q,ǐ�z��]s#{P��at�yt��v=N����ku��l�W�C����	�"f�N%MT�P��&~�V�'{a7O����3������+߭# ~��[Yϊ�Bo0��PM�QK:0|p��c3 �D�II��\��s��2�/�W�c�Rxo(�$4�A�s<vx�Gz/��_�-/]ZVV����oHl+�C�~[�r��>1�S:R�G��1@�@�7��p�/%�z���ӥ"�Ș��d���ݵ���.�x�l[������D���%C=ٓu��ʁ���+~����+�4�$J�䛲���MpӍ��:|Xʿ�t)�0�:M����l9���-��sW�����V�c@K����RX;�d���KɟvBs �`�.��8 n�@���ZyT�J�-�P=�/ӿ6�0Y�球aݻ�5�=��AD��?��ݟ�i<�_TNo~���tB�}"K�����]�!)��B�,�(�n�5�}�Ζ`çx$��4��� �/@_�C|Q`]a�ҋ��{m;��]
��|��hI9Yo��E�����m^�r�+WO�|����Ǜ��=_pl>��@�?�fv����S���Y>�T>��+h�փ$�uYҔ�T�+~�3)ǹޒ�I���>P��B�j"��Z��næ�S�_��t� `5�"���V� �#b/��{�P7�A�,��P��z�*kbA��28�ok�YT��Ъ�a�z�o�/pcف��Á! ����������u���Q����g�?$�7��0b��ΫƦ[�?�I �>[K>��֪w��%S��%ܻ8�������&�q����X-�w�2U���`���n�����Җ8��R}v���uK���`�a5c���?Jb���@��O������v@l8�r�"  ��P�EQ�81!�+�>�l���"e�����A�z�G��:ݧ�P�c�y���zǇ���þ�5xE,�3Q����A7��o�������;P��7iz=lG���ޝ��,m!�C�^|2��r�� !��e@���m��U<0���m�ªb�D�K�����֠�ۀ���/'��t?���d�G[w��>K�bN�y�*lG�@��eCC�Aʄ���ϡ*�pQu��>*wU�(����Q0x ����a�Ԛ���X�q�"����,XRi7'$���`!��@��]��TKeIA��`9��r���"�We�h�]�T?z��X:���v�cI�<\ё1�M#�8�$�t��Ǒ��^�xz�s��cqE�{{u�a~�	�fK�R�L#o�@�o���'F&��3���v/��-���۝=�%���S;�>7����OV�P���5/��SȮҜ`���:-x9�@�^�x�2��2� hGi�Z ��l�v�2���	�z����?w��#�ۣ���9��+����P4謊3���ߤ�ۜ�'~���%_�B#�N'ҀN>�������b&�Y`d�8��9-�o�v����j����(�Ex�R��p	��Pϒ,L�B;k���0���iSx�<�S���C-^��\T�]��0) �ۗZ�e=˰+�����b>QϞ�Pщv/3��j���dN�x���ux��ǵ:PK�S1>���I�n��_k���o�����w�ѱ���:�b���,�����[���8x�vƭn:h(G(��:}���8X���T�ہ�@�S���̍�7(nN���r^Z��bN�5�?U(��ҋ�A{�[�7�a��?�n�6(e���c+4z���Ta�[]]͇|t_QrP&\��S��;mr}�u�I(�W������I��A@k͕_�mA�f FG�Y�H�K�=�E��C���bٺ"S��!I�<mՄ+g��819�������R�ա0	n��ovK����ͅ��"��1�{�F�%:�xg� °��eW�M^!M߄��?b#����zRDSϞ�ED�NOH���D+��{�?��Wۯ�\��%��2+�0l0����p�߀�S�v:�M���~q:���n����[����ھ,�'�N,{\�s����)�B�L%��-/1:K�&�d/�us�E59� �W;�;E��FD���=������U}�)a��pR���_�����Ş��B�Bf�y�0��4`~@9��0b���̂Kv�8��-3��3K�Q8��pS���歴UC}GeOe�.�Fk�o_ϝa��-�~[�����\�m_�w�,���@S���.�P�":�:!��L����U��Nw����&Ɓ�jX�uTB�#�(*ml�	̄�T��VG a�g� ���{j$�Ӏi���S�� ��x��߅:ح�}c��1V���E��v�w�Ɂ���1�L�P�ϣ��GӣQ�� �th#oVӡ��"��<[��^`��g}�/�a�_�y9��=E��t�#Po+�ZC�tP|���U��);�H���_}X9�>2��J�:�ͬb;�HN?�%J��KbW��s�ֽ�UQסZ�R�����V�)�Ѱ�xuQa��|�Y�V˥E��9�b��)<�O��$�@�bL����������&.�Y�t(U}�� ��̲� ��'��7�����S�#	A�
j�a����	-��s�;$g�3�M����֠S��w�X���y:(�~��}�t�BT�v璡����³_�(�;���҅��I-M� Yh |�4г�)�f��5�v�E�J��~�p�;��PblD`�k�Xl&sQ�yO��~'�.گ[ � R��v��}�P8x�O�ao ���	�]�I�=��l��yU��=�q�!��'�w�cH�B=62�H7J�[��2�A���^8Xl��4����ɣ�"�,���䍮t��}��) ���L
Ƶ���ߠ�Cx�l	3�ߕ���'^��	の�
1TY���Ǿ't	�H���Z{�|cUF&Ӂ����!M��z�ik�	۩�wbY�b&��.iC��B#!0�N���c����?��3�n-u����î/�=��zJ)8ue���փ�ޛoXf�	۾գ�/^�)����M����O�P�3�*�]j��~�Q������~�(X�UX�zi
T�V,b���DagC+����@q%��z�p�AU,qE�?�}�M���/��8���/��x\�~��n�0�
����+U�,g��v�c��-V��uYDA10>b#bW��{� టs㶒3�����#�֛��[n��W��R����V��AMK�S��rR��^��?��7z��2�.טl ��sy�g�k�6%GI���`a��ph�v�D]y�AQ^�ڔI��!�7 ���^��3�,h���D(���0�:����� AQw����nR; �gÎ�^>ģ�����Gԅ2ɡQ>�2�������AnL�#H#�C0�
KY�M�&�;t��]��.;�L�1�b�Q���~�a����w�Br�!��l�kT2ϒ�����Š�ox�X�02=�BЉ��.��H�pM�T����*QɎxd�n��}
� ��P�bʾ\:TL(���,����(X�%�Ǧp�:�;Q��A���HgZ¾
L+��%-;��K�u�ȏ�c��x��cY<�e�z>�qNC��^����`Ș(�:}f,<�1�sl���сԄ
����n�K���ް��X���*:�)�4j!�ЩP�P`LL3��+�F������w����osδ���5`I\	 ��o��Dѡ_{acg��8�����
'j�.�Hm�1կ$[�O� "�D�����n_���䇴cg=3i��DM�Z �|�ZKɊF� �
���]�!:7�{��9�t�ɯ)�׀������E~^e	P��H������G�unp�fޭ�����n����D�U�����eQ�^	���J/�#]�󣈓����Q9^��F70��"�8�&q�%̯�ɠRx�X��_��LD�;kEmj��I (���q�6TOwD�3`�oo�G�;6���M.��<��=��@ ��q��~�o��Z�u����۰q���F+����FR��k	o}�F��>y�U�y2ۓ�1���θ�M��j[_,��\%�E�D�tˎѼ�L�=�h��L���k�M�1;�ʎ|�.'$���B���5#t�U�sv�h����h�mj�FdEݸ�><JC�N��
Q��xq��P��"�cj�bb�f�=In��2�|�U{�s���]�����omwrF�x�t�Z��t�-��R~@��J�H#ȼÝ�p�<-t���6��)`z��v���=N�@�zd�=�@#���ȣ{�2o��*����X�UY^��!��?k\)a�1���*� /��Y-R����a�p�J�a���j��Vt�������`�+�ե�Vj2Xiz�����ݨbV�����[8?Mks(d�v��
	ޏ!���M�P���T���� 
0�R�IN��I��	�b� Mo��\`�>�F>#/�XU�]H��k&�~{�l涖�P�Ǫ вQm�8 �PF*�Cs���竡�s)A��ݳ�h�����s�r�B��9�'_^�>�#��hi|2���#��������t햑����8u"�{����tzWi~�c����c�_|�EiR�}� ��J���+f��ں빤����,Uls�p��C3-f{�?��(�����]q<�B�����n������!L��% X��1fUJ����PЛ���L]�������xџ� �(�|�|+��q)��{x��+]�U�t7.��	�r*{f�'YCi"A��D>�g*n�p�\[]�-m��Zx���Wĭ�����?�j��'G�<��>��L��k����[��b/�|,��H)��8�0v�"E�@�:��αDы�<�p��۷8UƼ��[\J>sx鼅&�8\�ѧ�̻�u�W8�G�p".K�uv�	h����Qx�F����_W;���%���?*�?�ai�	���L"--�����"-C�h݋����9!���I����-V�NFpk�����5�b���y�InkJ:�Na�r�GD܆�V��s���5�+1LI�;�[�ǤMf���w��D�_d�iob�ӆ���KV��T��T�+s���<5��k|��:g< U{�Y�<͠�[��b��\�9�T�޳f�'�j��~H$zw�,B=�5X����5M��9ƃz�<�Ӫ�f��߶��WZ�|�8k���Ky1��[�<����O"h���\z���*��y�ޯ{���!�G�7=B�v,ǰgI5�|�(�42��K�=s���)L88f�^�`@@+XE8`������bi�U�{ѩkև叽݂����V�@80?{�O@¥��������g���},k���(O��=��7>���kR|4V���v��W'u<	�
9���z|�S�a����ص��m�UF�FXW�}zD���v}t�fc�������<25�߻?��2����ϗ3�#�k6o� ƪ?��.߳����R�<ׇ���*��#�ȡ�bU�)v^#d5-'����ק�qp5��\�k��!+�(s��AY)��g k�.c�sCt���$A@�u���v�ȣ���g��[V.I.�Fe��Y�̥���6��H���9�qqd��gBx;�ٔ�m诨�qw�}�)2�Ðgݧ��Tj[�|���h��H��$y�Έlbor�w�x�Zlv�æ���pH����NK,�u8�5� |W�r<� ���/�eߛ��g��$2�4*<Tl۴G����ΛCiKF�U�8�b=�fkm��U��.���#�jW�'܌�ZJ���뢏�n.lg�i7=��,h&=G�k���C�*kn�
4�@�R���ܫ��h�NJQ'SVS(�U���o�T)_-�o/�x���F���3��c$���6z�3hS�k��H�L�9U�+u�8� ����|�$f�����=�.~�����
�i�2H���6�Jb�n��ȤeFr���*�N�Ft\�2u'���c��~���Q���9ݍJ� �I)��!)�[�%�C���
���tIw���y�<����^��}��}�u����R�L�떓Ō���a�)%�:@��8!#(���G�b�DN�/uD�����$	�B���6X!��a��`@��6I�0r��v��t��T���3[TW�u7Aqޕ6�����,u"��D�Ԅ.�q-�/������8��?��z���^�=_&��:Y�����~@����}���==g�=���,*�[���5�H+H��|,�S�8���3D���vh��gA�[V�����(����y����>�:h���K��h�!��#����5$���ݯ�
�����/��(	�+�u��pb�o��^�X"����.~�l�;"�sR�J������p:G���j�D|F`�"S�l��+xO�`�>�_��O1�	]�B}�U��d�U2����{]~E��N�� �e/s���*S7�?ڦb/�unXo��r��k�V���+��~9O��P�w;�'�������p��8�%�$4|��K:C={�@9���{��a��O�&=w�L:}C����
W��w�qwW�B֧�2��n�>��uϯ����RI��,�g��f��$�"�
Q��Ð�,K�(j�4��+}��WY�����i���撪J��{����Xfz��(չ�ȳi�p(�kjϒ<~d"i=6w�Q�7�
�+"���|PN�������^|p���mM�+P@N����~���]���<n'P�On5�n���qZ"��'��m��5��(�-� ��9H�BIѲ��G^/�d�	��#������$㌥ִGb:�Ōx�Fq���������@H���f���Duh�jܹFօo4���}�}7�}ޥA�������>K�$�ƹh���j�/J����Ka7�ѧ|�1�Ą�!@S�1�ə����d���owߟ�*�5�
Yf.P��OL,�����jI����D8C�>~�ĕ�D2��+K�r5V�m6o�[H�/��r�;�l�6^��� ��O8�H�	9���{Q��ν5����>֣&�n�,)��p�Ɓ���L��K��#�6ħ
�ɗ�ː��d@��!�R	����^X��R�Rߡ�*|@!�e�r��?0��'���e|}n�4*� �z�3�y������s��6��<[g`�w"�5�a�_ -��2��$�G�g��EP�~M�̲��sY��O1����B�S�l ��̡�?M6ҏu�oם�R�')G���œPP�"e�:���*,��}�vm�r>y+0a�͐{���O1�vH�^Y�f����N�w��_IL*���Ҡ)��	�ҭ y7��f9��6�CZ�C"?mq��nas�1���Z��gP�Q-獼ʌI�2��RnTjk���?�B<����o�X�����3�%��v����V�B�y_Y��"2��S�m	
}��j�z�EX]��{XԐmK$�qW�G�n"
��t��̋�}u����V���L��J�mB�n�4�}����?@����Z��zɓ�$��; �ǻ�I��\k3�R�su�惝$�:��>itc�T��~����Y8�ǁ(+8��ut�U��ߒ����72��q�dƅ��^�Upy�z�/a�A�?GϗӠ��hY��o2�&[|$��K����4,/�J��1N:�D�ɓ6�2�l�$:lh��`�._��-�θ\�Ml�N�s���($]�)��g����z����k�a�c�D�O�q��ZS��E�{c�'j�h�!˂�����r����uOjizY���+1r��'�w��������	YX��E�:�vv��??��_�/M�_pOآf���;�O↔v��ء{�@������2U�s�+$�v���뮜��/	�QO�[��>ƿ���4�:&�c�ן&D��҈}J����G/��Qi���=�-��v�b2�Vi��K�5�"h��� `���
id{��9;�\˵����0����W��=�H��&4���Ғs�M�}4n�N|�����O�B��,Ug��8�v �r7�1�0/��,2��w=��?mY�:T�$���'�	��}���v;�p�'���W��� ��_��-�z��s`u�~~���v��T�|/�}Kē�ؓ���^���1��u�#�M��c+>�c�Fy=k��\g�1��I��A��O�[�;A^�K&�z ��^���@]Z���{\��헴�(��8]��/y�/y9���x���'�+T!��:pFji*x;f��	�ځ��l޼]����%�h����/8���:�|8?��V�+ #�J�%F Y -?*Q�'��䅧�@�{�:�s��ax���xT
Ps��]��{�)��Ѩ����@��wֶ���i�D���}!R�ͯ��⤸�7x���e��B��H�_����΂� ���@_���|js�ɳ5w |+�t��K�~r����.��ڭ=ۭ��j�X0LԷ`�Y^_�A�,�M��Au���`��޳G3��M��˯g�G�gxIW�RxOtSJ�d�?~܁�����z6�L���ઓ�\G�3E =#��i$��,�<��
nsE��ʫ=��+8D0��[@m.
���ğ�08a�G��x�X��P*-��J1xn߻�(��D��C�)f�5��4�cG��A��掖ma� j|U��]B�|��N:��ý���/8���2�޸c6�o�B?\�⩽ZC��n!�Sz���v�w�o��87����/����W���S)���ޝ�ȃ�]1镍�@F�����9~��N��~H�!��(���U�g�)Ak�,���I��8s�c�=G3NDUy�2%��#~_n"�\��=���A���y�h/���<�v��)��]jҦ�
s=TW��̙3�3��������3���Wėi��@��� Z���ԩ�D��,d[ܶD���7�W�>�������_��?����enz��A���L�;�QP�H0:Wrv�|�u����/y ����a�n�~�+�㜰
�*ʹ���g˨W��̤Pvq�B׹֫Ƶ�5�?s�T�I���dN�vq {��n:p@���P.�ɞ���tsy0�5.]�jC-Q����e��F���_N�'�"!n����|�>Z,��q4,c�T14�?m�����"�}��i�XJ�qv���՜Hu ���/�p<�D�bLot�<�F��o�
�! ���/�g����ajJkU1W��K�s�QAF��Lv��]�D�O�k�i�������dZ��n`eaEj7�(��X���
_es�bi <&nR@�͜/��i"�	�@�h��~�e?�6*��g�*'����8�-s�8+�a%����JQ�oƯ�d{eܙ�I���V�uNZ�{�����}Ń}�[y,�&2�@��-�\a��F��,��yʸK}pq�����L�{���w�ޭ`,�r��,��u��^��{�r��u�.�DEQ���r���Q8pIe%2��"*1Q���b�_è^�p<�R�ӫb�3��'�<�Ӏ>��܅O?��):�YT��L�m5�f=�T�
���s�&������j�z������alˢ��J���O0�˨���~:��T~�����h A����n�o�Pͽ�5߄��/��o^�֎�`-0D�LR�
N��8I���KV�?�Yj��JD.�)�[���)A��/��7
��3��Ơ.�N�z��;�!�|�jo�9�5X�q������c�щJs�2-�
�.�c[*6	�Ƴ�E1��4��1"#�rløaw�y�Յ�4�	����n(���\��x�a���KNQ��8N�{ L+�9��0���+t�i,�6G22=���%�i!*/ƒ�Ø���a�A6 �tO��e��HG��Ab�(~��8��V�G�5��fD�x�]�{���#�7o��� 
� b�(�A�/بPFe�7��X���0�Đ�	GtU&�'��k����W�1��O���v���V�'��W�[?�gL{��{�a�%�h�Ff�bE�Bc-�@���ܖm�S)���\7�;�}=�X^~�b�-=�����CϨ7S��^k���������uH)]���èxWS��
���T�꺴�z��w#�&�dm0��� ���œ�lONx��A�<���꤮�y>�Ğ�O-+ͳ![sH���x�E��V}N[�u�����S�*׹D�|� =��t/��=�����m�%� ��}\\��<|�� �!�� b{��'1߸��++��P�ϒ�/y�W8LgӲ��&St��c�q�����$�[m���Lk!j@4-aNT�jE$����d�����2f��c�,���7�s���8�r!k�k~D�����D8���O�w�
u�U�Hi�/�8�D~����t&?����t�z�Ħ��Ъ��$.��g�pD��wI4n�]��L�f�$�� �V�?!f����o���Yz��9� 冈��py�@j���$��HO�U�)��u�ܕw,$��z"AR����\/X�!Tk}�p'`�c}�b����<d���z�yr�!��B&����}e����f%�4���u��j{
R�̂�%r����>�GTbFq�)�xX?��}��\���}n-�fN��ɌHmEJR�vel��^�j����\���}���Bg�QCg��N���ޗ����7A�Q�2`�2�c�9�\�/�.������m|��]��$L�Յ�_Mꬄj�V*���B�����'��|
���"�����Xo����q[�Ax��o�_%~�n�G~(d�$��L�+�Ui�"�G�������w���Jw��~��&�BD��eU�Yvd`�ho
;!Z՞��2n�k(�}��jB)-��\�	�	R���/O�CI�������I��]��&��ǁ�?���	"�����+�����
�x��$�S�[VT���Q������� ��Ӂ?�B2��4]��)_%�X�"M�U�>Zp8�<��0�N�Cu�3���	Ӥ�&�@����N�E!OϮ`�{��R�ԙ�'�@�wp~����r�O�����I������g����fxe�a��ӡ�3����J��|�>�V|ĩA�1��B�~���cDW�]ƞ�{�a��\��w��&ô�,*N&�|ʫ�xHu��态�OH�*���_�|�7ʪ�U��z"Q�s͔x\D����H�=�&z������C����饩�赼��u�+�,�ݗ��X�V�z��~Zc��X>�ƌ�]������L��բ�B�ײpY�[��l3L��B�;�C�I�!��
0���N��Z�uގ�g���}��*��"@M�L�ػ�$y�i���£A�!�QO7HG�ڞ�V�>��"	������ױ��0;��Z��l!I�pG��Ä��qw���Xoo2ra��{����w��X��P��/�f�d�޶@ﴜ��ҫ�(���ߢ��Ǭ�4��(<\�A��[㷤LҲ���_�-"�H��TY�z�x�1��>ȗX�,�u�������ЂX�PN���7�{��܆���vg�\���s�*vqh�W����Z��֭4��璊�6i]��S���[H�u�>�ǱZ�Z���?l5i>ۆ;���n��$�L5@7܂'�䜔 Go6\��>|��,��YA������tM��PWS+;� �B86eW�\�:	|%AX��*4���K�j|b�(RFp�>k��x-4�[G/C����������z>N�gl�����V"�q��&޹��+~;�:��CĬQ�~ڭ7�y1-_e?Q��"����}��fhzT'{��d���2�D����t����CƊ���:1z��}*��@G�o�r��0�W|͔��f
rHkq���=s"�m����Ƅ�����(���S��g�l�Z��N���V��Ȣ��n�6�\�Ry�d�:�ŜxY�s��L�����[b�З��z�_|�G�.�F�ی?�~1���|�q	nw��EK<8��|/K�A�ŦR�E�3���rAe꣇�Ia�u)�o��������Kb_��ߗ�1�=<�p�|���!:������
XB�8�I�d��D���i$��/L�&��a���~"!�DE��nw��1�u�>T����qU����ԝ֋� �b{�<]«@U5���?�A&#�^�o��j/'��6빗䘒�1:fl!qd�Sӊ���MH��e�k��+2zR� � �r%�~APi�D:�T�;���M�/�U� ���er:4���h�+qx�����Bo���K[�^DFeڨ��/烒ڴ�*n��]@Z����k$-{�f���d��.�PY�*�&zb��׎��8�%��);��!'q�8"1������n�{�C9-�@9��d�I�������P5FO,�t��l0���-���Y�C�+�m�N}@]��W��:ƚ�A���k?���|����k���#CHT@Iˁ�N"�B�G�`Z��33���BEy��c�n�7W�����̠��F�����AG��c�OZ�>���O�k�oޖx�`�4_\x�]�G����±�n�1 ����ɱN�rw՟#��5e�5�0���
���A�o	���.to$�:�*�_v��Bfճ�xh�N?���8M1�5|�=��rҥl	0F�+�\)��0�.��D���~�&��/��*��.�s���Ă���<a��p�f�NJ�$����s,a	��+K��n���/I�� ���lW��~�-����ۺ����~S]k�n�3c��ń�E� {�e�E������^:�F�����f���0�⋁n~2���}iC�|�k4�t�5[b}�ߑ��%��`����UĐR� �l��_Ot"��������fH�U$->	=�7Jj<1��"CHI#G1��֖?-�_�g��H
�Kc2Ti��%HQ�:��0} n�����G�ŀ��}����*Q7D��]u��
��5o5��g�u�S�#��Ay ����!-~G!�
ς�i�����~�yH�%����sb�ɍ �n��=��E`i���p̉
�4f�؍�&���sH�4'�k!
����ѭ�����#2)�b�;�sB�EX��$u�VF�Y���J,�bK���v4n��t����j�O� W����0�t� %��]���s�եJŵ�o~����M,O��Z"��N¹�����4f4�#zj����r��凶��Y0�8{n�:z
Lfy�铅���i9�<�XKeB/�6�Z�7}C�<ti�mC��wOn̑��JZ+2��0���;p|I7�1��;蠹�rf;>�+r�	��m =|����kd�S@	���� �ڽ��BQ}&_�����Z�ybnLH�=x��ɣzW#���O;�5�����@t���ߜ\џ�RF� AeX{��<��Y���Pm��9��;i��N��b��"BZs�S���:����6�RP���~�A��`
���-��T�0\� ��6e]q�`c"�m�T��7Xw*�<r�Z�jLU�Р*3)1� ���6��t�&@G���Q)�b,=.�r����sv�8����xZ � 
�h�J,�:� NK��]~
n(0vN�	��I��ߴ���bQ��	N�'��-���ogV��s� ����R}jX9��uUM��B�#�v�E�U�!��eKq��;��(�p��n:��h,��	'g�MUP� �c-��x���X��N\{%Q�����x�B���R��ንa/h@q9����]���(�wȯz�Ę��Q �j� @���?�G�"�UWq�����J["�R4'��ʑ�PkZ��pJ��I�Rk��Z<��e5�w���w��|@�XN�"��	n�5�U@ɧ����@��RY�����.�����i$M�" ܞi>t/�����ww�J�ў�J�e��\�|��ޔ��ڸf�*�bDM��NM9��:oh_����i.*�<�`0X�#�YSIJ�o�������+�U䬈��L��P���QFɧ�w�D�����Wm� �R� ҩXLXt�bi�"AGE5 c�t��_�M���9���;ϕd�mƞ�i��?*0k~E��.���h��n�����E˹n� �����H&�BH�,��'�{���;ǉm�w��#0v�7�����io~�0}��3�|����U�1dXA23'���?dp�o�k��(BFe�;~�����\�[�t�w��r��;�)i�"��.�b8��~���/8`Vsӓ��U<c��#����#�m� �WK?d�1Q>&ԝ�1|���e�}a���ź�֯�+���0pY}��!��Ps�����,�1�*�םUQ����Л���WO�[��0��%B�"B��#5�������1bļB��7{�<dD�4��r�Hz��¸y�~.E���9L-d|К�lg;I�KF��J�h:��p�	<@-R��M6��ゥ^Ĥd�C�B����ϟƝ���*�6�$_ժ��}�&�Y�T%�2!G_���輖��n�N֥��R_�M�gz��Кz+����zi�kx���p�8�/R�+�N����X���j�T�&���򋯞�u�j�#��eof���1,���8�.��v�L-���3�W�qۖB(:,���r�T���\��B��2橎Ę<xaF��&�6 ��� 0:�'�����
�-��b��/�Y%�EO�ĲUBx���Z�7[|���*�n�}�F�Ɍ�`o�|��p�&,��ƗG�U�$���	I;��T*I��5�a�;Z��/�0��|󟼀�G�._�a�Ӓ`1�&jM;���Y�; 36�8�����Oo9��x�����P�Wr��W�0'�jDw���:ד����`��+���vh͇�RC��}���~&l�~�A/�u��G�0&��']�ޘ�� �]!�n-`�au�չ\���}�IF���� ���bLuջ�wsh��I�C?�M�z�2L��rՖ��ܖ�]dl�>aj%�Ǉ�m�2�S;&4a�&�X��W/��x�U�ߓ���!�@�V75	��|�Ar��V�>�%�:�K�hҎ91�x�=ᒋOkV��g�ԏ{\�]{ |�=>"�3��m��Ba&�`�oj��mM�dԟ�ħ��6N�̠����72��k&���왑~��
�Cx'У巨�,��׀��˿��Zs���;�$�H4�#��Q�j.$��c��c�(��Ur��(sL�t;���4F1yL�4~��_`�i�@u�{�N�kC��ܩow��Ն\��u6x.f��b`� �s>�N�֨{'�F5ZN��F�6tў`
�p� �"H@q1���u�{�9�_��!��;O��A�$� �����IK��GF�h=�m�w���5�r�!R3��Lܼ߸������^Dn���w$i��\R���y ��|6��"�N���U�|���	�x^U��G�$�?�L�mN��#��sC����M�;:� s�s��7/ϵ��xN4�����b^��Y9ٍx:�8�Ż����90-�]nN�y����SA�{�E�?܁��������0�}��߳����B���w�p�����6dLc����%ǖC�p�N%��.��^�W���X�!1�C�2��\���3'k@ξ�._S'q��c��c�7\�+*@�@�_J[���Ϙ�·D*wb�E��v0�\��6�m�,�a/��Yܩ���0v0���;{��_�Y���'#�eK���������:�p��Y��=cɵ��ToO?j,�<�@�M��8���q���I��������}OQgg��G�Q�kb������Z)���M{�j��� M�6̪��!$3�RW��]�G��N��6p��7�_�5��$_җ�(>���S�NI� pWM� �\�٤nȫN�X�e��ۊ�����qg�~�w�����~��'C��P���ON��Zv*�H�1�Dޞ�ey�e�]�qM���M5Nϊ���&|A����5��n���]�ҍ�����/4>-�#��}�E��D0;XGs�7��	�	��! ���t*�*(�,��$U@8����s��Y�!�L����4��tm�-�@\IA[�ER_�W��),?�3�ך�'זX0Ֆh.G��g��6I�o�%���'寊��$nY,{�"��=���[0�z���Af�fR	]��[cc)qP&�'��vR�c)T`NA���!�y �ٳ�������V�	 #�����Yg�oG@��f�E@�
Ʈ|���/�,�q���%���rp�>��ɒ�2_`�@,��}�齣��B5��	v&Σb ��ɑ�
sq��ؕ(q��������'��R���킑�>�A�r�o{�>�]��_�"��*�� �&
���V���8Yx"��
�oYC�UO��� Ou�A��&W,�#���^��!���f�7O>�:د)[���� �0I��O�Ӣ���lG����_j�n�=>ePXSZ�r�����ܨ������~���3��5�E,�1�܎dV[t0���ݵڃ���k�VH�%M�ڙ��m&yH5/xu-�r��#}�|�)�v�]�Jӂ�f~�r��g�i��V�m�</��D�([��O,%. ��]���+�����<𚁄�z=�f�:򣁥@5�&��]�GD����� b0�3��g�D���R������ik��r�f��!Q�sm+n��-K�	2�Sd|��z�.IЙ�uG�c6b�l%�y�`�����uVܿ٬�b����D�h�&Z�{����*��֗=�ʺ	{'��گ�3���h+|./��(g
� �+�0��(0}x��R�'�~�<toݵ��wM���1����SӶ�҇�a�qPƞ�j��d;��gЫ�*N9n㦑$��K"�_��ޕ�I����Y��� .z�j"���?�{�t���,:���4:�٘C�7� ٲ
x1�9�l�y�<��i��F��a�d��g.��"]�l��qw!;��%@pKKW���M�$迱��מ6X{��F���E����}r�jWLl�1�f���(�E��LH���ħ�O�O[[[�b�0s�E��J�w���{V#����������h8e�TrD�;n��¾�/��Mz�щ~C�
�Vz�L���*b��-�jD�!�}ҿ|����r���̋�	�TS�؆L����>XYe�o�h��@��˒����4-�C�v�F�v�$f���p�=�����0�AnM������ �r~��dð��W�K�
�Ҽ��RC,U��r#����HZ�OQg) ��K�xvi���w#�����?��ǿ���)��ŵˉ=�=KE�tZ�P�5�(F-���~�5a}2��B���@v���}����4;�9U��B���e��Aѯ� �O���NcO!a�����Єd���"���Β%j�T������}k&�~�z�9gN�(E}҃��~�ў|f�lzT|ڨA��1���%%t[�llU�L�"�6	�8�=��=���y򁏆�a_�Ά�`�/+wS��z��aӗߜ��X�L%͎2���]��YΗ:B����ZbM�)��4�da� `J��f�q�	'V�4�m˺N�E��d>��h�u�#P>��~2(���)X�/j�Nl�	ּ�;�s�9'����&dR GB� �Z��� *L��~��vXO���)gAV� ��.|w�]��S���J/��l
I���?�c��K��.��G5 H�$H��c���ŉ��R�&�	�8r�9�ܕB@��}�i��FǙ4�
�o��j�{m~1ܞ�7hm��6�������	�[d�2����A�i�сWL��Uo,o��rE5�0U=��cI�q)j�[w��R��9,h嫌���2��2��&9S:!�y&Y�?��|VjҊc��^:;�}e��W�\���E]��v�?|�$S�^q�0M��7�ijL��v2Nқ�(Q�<�T>a-���E���㿿J,@f�oaJM��*p+W"�"z�¡#���cô����I��ct>n�D������x��R�6#�|d�Ql��_Ƈ����臨}��	JdD�|H�?�Xg�F����B�O�{�j���y�U�������ϙ�}��C��H!���z�p�~6ڴ��l��uA��3���Au�R/�Z�m-#mf-��ˍuF�����'IE��M���rk�R�_ph��F��[��S*8G�ݸ�X݅O��9�"gE����]yk�4k��s��Ʌ]8ȃg-Y������V�&�֞���jY"�f��mA��T��?�Wl)mU��ST�X�(��V�l���7g��ҔS�(6�C-��4[����������w��:5��r�<����� �`jxv��@E�f�_$g# Rs ��M����> ǣ��H���hc|_����ly�0u{� b������4ه��Q ����ɉ�o�J�JB��/�?�|�(XKu��'(�~��b�^E�d�Bvz��� 
޺9}=�9��ok=���l��:h�R��}�6t��lԵ���L���Y6�JWX 
w�r�f�T���B�:���y�]�%���#��g�Q��}��f>�Z/ί�;���2O�c�E�E_�^Ϯ��~l���� �?��|�tAciUoI�x;quuZp04�����̰���u Oٍ	�,���@�@{�o&�����p�S�7;�|��2�=	g�4�7�Ϋ���|"VM��UvA?Y�f|�C>-~�i䂿z$&����Ƙ����,^A��2���Ć!�94�t޶";O�/!]m���y����L>�P���A�E����Nޞn��S	c`m���������(�ϯz��K�lT̽�T˃6|֗�#_�ƅ��KCwX��Ew��Dd�͈��y�)�N��N��j�����Q.eٰ�F������`����JE��*Ž�N
Ei59�Ɠ�<,��i�^�}��z�r�|���-�r���o�'S1�'�I�×L��Љ-�~����|P���7I���i���
_�"�D?g�e����q��ߟ�>�*��dˊ=��L�
t�n����]ٺ;v�y���R�ǥUxp���r��3�R���`B��`�zĽ��)����6!{}4?-P"(Zp��n@K��7}?NI���J��\�>�C��Z^�# �7F@b6�4R}�^9�h�j�O� / �G\5�qu�?ʥb��|i!b�དྷ��;�������'���؃�K3��mU���y��#Z���]���Ӡ�S?�}�;<Η��B���b�#OM���Y�X���Hn���"��''�����4]��[��1�ڛ~����E>�7�P����ǦEN�Dįb�z9~'׬k�{��-���+�	y��_YLջ�����`~����º�o��V|���T��;��"�ـU�l[����=���,��	Hh���!80�BR������3��u	Էv]�~��rU}/��y^|��&I!�oL��/�m�h{�3�#H��0f|s�̘���hO&��lh�'h��&O� ��I�l4:`���8����-���4��f^��S��0�P������x���@λӋ������&i�E�I�UG�)f�М�_f��$�T��_ډ�r(X����1�1ڵ��1�΢��>�_t}�-"�)A64���e�P�C��nq�M�0lu6	��P�̰	I=��J�Ā�ěv��<B�����Q���w݋��`�b��F�'t96�^+ߑ�WJz���!� %�]?���j|-���R@Km�J�F�Y�x�`��C�.͠"D8�J�ۻb��6Tǅ�� 1�����4;U�l�+&h���x'�7���2A��q�_�OD]�B��&��a:Ƈ/v��¢��~˲v/�+7'k���w��n}�E7W٪X7s� �E�Φ58`}P��dʽ�jT5=x��` \�MR��IJW�2�U�7B.�|��[��0I�ϱ�F1��4�4ft ������G��A�Z#���-̿��D_����ƋuLVl�Ю�]�n	�������>\�ח S(s邇:ϵ^U)�8�������9�ֿͧ�M��:%��4i��f6#a�:QJ�j�ƃ�j��bD�Z�c��&p!'mz�X��i:"��� �3MdC�F�	�O��;�\���x66Dh|ڥ @�Ae��ī���bm�|IJ����W�%8�?`@g�42��]� '{它� �=���qƊ��Kؘ`���	�	9[��Q8�Ҍ�ly��W{;O)���|x���<�]Ϗ��ń����*	I�!�������j��Z�E�ٍZ���E������퐤��ܹ'Y���� ��ơ;?��z�V�{�Ů|���A�;U�~(<},��ٞ�b�utYf\�:s�~��M��1�
��PoX|)���9���D�##&�^U%=_�ڳ�?����q�%� �9�%A��7��,ݍz�fYɺg�W�q*%|ԩ<`����<'�<B �=�w���*�`Χ��T��I�[�ϝ.��?yq5F?xM��9$��p�Ρ�zT���U����f}f?�!���͸��Vw��L6�z�_|�N���}��ᣣ�.�o3�AmT�^7K��R�#�X#Ώ6ogO�\o}	�2ïl��(>��r�B;�!�4�ND�6M�gc�Z���y0A^��kF*����md��!�F��;e�/&��2ks�LJ�i�g�*e���,֨�<�:Z�� b���ű���=�Դ����U�zLL�83�ծ�QB+���ab��x�]��|���?�/���V���`ߛģ��rudvv}��0U�Jf�I%uH�Ք�h�D�(����iR�lY4�l�Y��A�5+���P��7��rꚵ_%���ź�KӍ^"���h9O���>���1���)��D�� �:�����5�NHxWT�p"��(�y2���޵r+���}��o��*��*pͳX	�b�rd��]#p�29�������$�����܌��/K��!Wj�W�I�V�?�tz��˂	\/Jg�K��ܷͿλ���l��ވd�RV!�x�����/�(cF�F��FV��J{ߨT����:���>w��щe�G2svG%�!�
���"2@͋\3�)PSq2@T�I!���6����"�دD�1�"Ya��� ���+,����`
(ٕA�P{�y�izwyOE�������+]&��y��+o�"�1R=����=��#���1��i�z�x�B2A���x�=��^�6u8�g��<�ZWo8�K4T�:�3:��,o.bE��-~���Æ����m{l$�1�!㛒��?���ă8��fD�}]�To�4A��ݧþ�~��|wP&
�����<#AZ#խ%cM��j��>�F,
}�+��]xI���; �̈́E�~u*��&� �9z�u_܊��'$����G"�X���ɂ밧�X��B����	�4���i���F��v�@Ӆ�8p-:�xq�~�[d�X|+�b��|�2�s+�6-��%�iB�|�{�"Ǳp�Z�)��S��@{���NHۅ�`hT���QaKd�3����.aҎ*.Q����8M�2}�U$1������9��v+�#�7C2�L*�:"1�/S�B cm-*f:�v�)F0%��j�#��������R��UTZ}��v�uӽǵ��A�}�a<�x���Z��gXl���g��x�EZ���vW�I�	#�ҙ�Zw}�LB���������>��]��K����;i�1쩣�Ґ�!�"M��s�(L¡����3Q!�_Q�	�"��k� ���Ӽ:�mx���l�}Q������zv��W����Y�dy_�鳕����4�%�3hoE�<����!���9w��D��\@���}-�й0,���+s�E�:����<�`���c�[�4�mZ/���gT�;��\%��O�gr���x�e�>Ɲ&��=X���|3��|�t	�/��v�#��ޣV�~�]�=|��bͥ�qv��=6H���s���m~�(0���-�k̝���`I��-�Gɏ :��{<Uc�Gk0���r,��!�b�g����[���M`�x�b�Y��^�b]k�ٍh�/�a���f����B�O�[�mD|x$pfM�7�폿���Ǝ�D�9��@��(���%fN�j�IX�"K3|*���G�l~z��p�1����V��@voPe=a�u$[��/��䭶t��܋�hV HR����
�*u�>��bQ[�`?m��쒇C��x�qXޠ�q"H�Tu��!�y��&�V3�D����I�����Á�?d7�8�,8<v2���4ފ���D�F�S� ֿ� h�ٯ��*�d~�R��4c{�w��'��vӤ	�Ȼ���86������J�a���O6m���3%��]�C3e��n�L�qZ`b�T�[B럥z�Y�<>p�uWM�����XW'7	��4�|�w	�r ���bs�l�?99���+�SS��<�e|H���=yܳ:�ߢ�Ew�qh����T����H���Сi��_ƭ�·p��l�O�����Z�{�U_�t���15�F#]�H��J��FD �ҡ�0R@b�t+HH#�"����y�����v8�����뺯�N���J�i�BJ�G�"��&�y���]-ʈ�%D0�������:�w��$~�Q7x���hV9!��[�p`ãC�I��0�_�9����c�炙\��9�P�I��a�����(��0lrq��\a�듻�
4��mo0���3+ L������������1�Y�"��]�}q�X�h���T����}�.�B���Y.�<J�E�Θg�����Q����`T��
��ӽ	/ԫ����h�g�H�c}=��l�H����ޔ�ˇ8p�
2�����g.��Z| j��_B�Q�H՚E��w1P}	��D�H�}��6�-�f�`���oև� �t�d��s.p���!�}ϋ��S��Q'.���������ڋ��rJ����J�p3��
?�E�GO>���� ��{����t(��CI� �y�V��å��k���6�kk��>R��֨_{�?�]"B�L�#�9�;�<;2k�N�N�beJ&�ww��@>�4z�$��[U�+�*���a�y�ps8��M�r>�Vad���F�f��{����UDY���)I�#&}5w���E_�$�8L�s9"E5y3f<n�&G���o����~F[=�c|�9�ա�@�XR�'�<5D	*��F�:>��Y{?��rǀ�ϱ"�I��BP0�u�6�?�������7ֲ�������Pr��L�u0U|c���_�ޞΘ�����x�c'ϳ=��xH_�a F���p��wd�ꁜ��t���U��Ƈ�+��VG'\���05��-)ӯ/%�"Ud,Z	ﶄ��l0-z�.ĀE�d�p�&����&��?�0;���=~��>�9�n#i��eÿ����$�4jU�?K��BU�^£�_�i�A�S�!VWA5L�y�5�JM��,]�'o�4
��=�L���\���a��3�s��W��*bIBj�&y�S�]��\�.���(�;�3V=ٲ썢�:��	}a�9��юḿ��%��7c���Bn',���B_��٣J�kN��~"8���ɇϋ�.��H���A �O6���c"xD�1��ֱ��0�zMZ����3m��Eؚ��ґ"̃p�L�e�ZK��/M�x��s��r#V�EbS�Y��_�ӡZ��A-���;��"�P�"����L켝�;3�j�3�;�!�2��uv$��|r3ߔ�K�IV�X�R4�5&P�����n{}:JH���9�^9`rF��k�� ��/�"V�=	��/�,��|��������{��+v�;)I��X�{��8����2�ങbf����������#�����)�]f��<� B�=V>��=qRa���3��
��V'V��h�t���DpWs	J�* ZL����]�q�0��݂a"^?�p��:���V{��MFrdf���1q��:��4���B�З-��ֈp�<�$��r�uv��W�}��4oAD��� �?�L^n�@�é�2 7@>!��#Bw��� h^B\���Awf���5P7͟����B�+��
q9��9>	������̵�U�e	6����ck�ƕ�Gw)��M.gN�F��.Bx Nak���M��,��@���#y/�k.1D����z�nbD:�֯o� >�4Ɍ��F*F��K��!��-g��\��>r�7�	�j<��43�_Cw�t�!��٤!��@�p*��+��KR�e�l�w�J� �y����?	�나����.!���b�������I�f��]�� �;;�4	���r>��%�J�{�J�o����p���x
4q���y�z�0�CvU���~y�'I����$Vw#P��� ��V�V�TJ�q-���Pj�#x����ԇx��{3�wS�X��(,��i"�>��M|k��ſt�&� �0i���{z `m�&� %���f1<��ic��rE�����Ι'G����Y���� K#H���GS���\�=���܆�<�#h��IF�N�iFaQo�s!���)ie������g]Ag¼��Ӯ³�+��:��p��a�oI4b�	�s��^E��x"���a�t�HW,F�^�#������4au��|;�U���(�֝�����\��3[o��訟c���MW�J�m2Q�Dh�6��!����[+n���] �?�q�k��SzǄ T(,:�Ԥ���`�;�d#{�C�QWm>~KHo@��i�hP���BD���Y�:����B���D:�&a|��qf�w!�������f"Zi��07��<^{L�|�������& �Q�+p���sP��ԕ��x��~|��a�����A�ϲ�x�Opa�ƺMV�F=�8��ӝ���7���z�-.��܊Cag�������+R��L���΂w�B�3��l5�ժ�I�"-<��]��~�5�p�v{���@��à�[��V�?��X��P�S"P����0܌Q����y*�ޜ��s�jI�dbH�%����do���:�e���H����3f��$� �.��?H�ve$N�~��/N�	�wV�_v�OV)0������vQ�����吮v����|�'ݪ��WV�`*�MƪR���z;���� >�_��)h�Z����g���4Yy����5rek��{�
)ԓz���؅$�����ܑ�R��,"*�ԡ�H��.���{�b�-�t�{ҍ�B��v
�Hn	5���\�C����� ���+�{?').|b/�\p?Y�E�8E51����0�ٽ�Ţ�Q���1�R���kp���.]Vw������ߑw�'�q�[�ڄ�I��;[߾�{�	�¶R_�
.��_���xL~�}"���1���,��Ҙ�j� Bs�����W��D����-o��$������zLf��}q��eH|��
4*����&��4q8�#P��<N�=�'�k�p��5,/�٥�1=��awI�2�H�^{gH �{�{�P�>���i�X�X�ݻl�)s���$�f�5��g�?E*R����b�lU�t��CD��z�R�����c��	&�{Y�~PȖ�Ì|����W(��ؤ`fPg��U�>+c�1A!Kʮ5;cb\oC� cʛ�^"Jܷ*}��@h��B<D��&�@ ��������)J����.1��;�?\`y��£e�[��U��c!��Y]O�67��\|O�#^P���'�p�ps&�#�T�(ǲ�v� s��Q�nQu�t��*��� V��X1�_���N��U�zM�~���f/i1��Kz�s��˨x�A��Uz���WQ�,3���F��,�욹�I-�Y���W8uj���Zv�\��4I�ߢ�E|��M��#W����Wm����c���z�$�Z�H�³Qu��_�B�j�`����ߝ��k��2�����+�� xVZ����H��*0W=�n�Z�G��Z�b}Q�?d�@4�qJ�CFD�Y�(>�r��D_w�'�_b:e�62׽#ch��W�"�J�J��ޡ6E[��'��|�W����ן "s�m�z���q�M#���3f9�����471n�����p��A��$���g�dH �WGo�]�)$FRD�v�v.A쎢���	~V��B��`f�e���m�,޹�&�с��k�~Zym�ʵ{n����^�Mb	�������̛5���g��
��N�0\���0�~|�'K�XV���(PfБ����[���ʅK]�}8�/�T�a���p�������)ez�1�Fo��f&}��������P �T�M�'���^��|r�?�������X�����t����0$x��==�Wd)�����Е�W�'��|���!$��]��҄u�&�<Fr���6�!b��%6dur�o,�AJLD��H�#?:U���L���3ˇ��*$�����"��}Rsۊz3R�Vl�UD_.�+���?��!L@���Yt��e~���#�ȏ��c���rz����»jSӌxĂ��+��=sη��{�hy�7��ڜ2O�+�ףYu�{�����g����h�U߇��On��M�lOn�	���_��L��Ng��+tu&VS���Sn����H(IƂ�Z3�����UG|u5�ϒ����Ĕ��#�����\�qX.��������g���޴�~u|n»`��13�֫A�}0�x�D{[�a��t�f��)p�!��n�>�q`���߆O�#k/R�̤@� Gk\�>���j��ޑ�U�-,�KI��Z}�~��d$K\G,�]6��yh�hQ�:9I����y�ye��g�����p�%qԑ��<�� B��fd>F_Y�^`�38G�!����*���¼Y��m'��xOI{{]C�魔��/Ї�uE���6��Ec%��
�=�i�	��heN�}� «�RΓ��n���!#�I��+_�B#����>���Ի���nx,�oV0�i����*�<�d7/���K*������n�-o:�ωߊ�-7���Ȓx>��^̑��$
k:qG��(҉�gӞ��ڬ���MϘ���{o��y.�<�F���Uh���C����כ��Cf�d���<��I5�x&��>�"�A��������I��։޴O�&�#ٕ���{1~yAJ,����^�%���$��pD�@���ơ�m�fz���jO����$���굲E�~�QEb��"��;���N2���*�~�קg�k:G	�	� ���۸�E����h����䍢x���e����=&��QJ��o�k[P �.v�C�ήR�(�X��J��X��x��#�p�#hܚ3��" �V���*T ��$7�@?�j���Y����p�ݴ�}0�u��aD�>����I�ˁ�^Au��SRD�-�!e�e��~ǵ3�\a���_������}ɶ����*|$��6��_�2Kn���q�/�ٝ�[`��dZ�e�D���|��N��7H�3+e۹�����t�#�r�xm��<��Ly3��BϾ�J�w�Ρ�ɋ;���ύUp��Τ>��--\����b���3	icF��I�Rx�4;Efٽ�ĒX�xL�s^�u:�z�R���-(P���y�*�؄�0bN�-,��=�N��ձ���Çl�8�=p���S���_�ڍx�����dKޛot���t�$V�\C��),3�Rb\_{U%�`0�r�5y߸�'�4k	z��p�n��@�h͋H`p�G��zoq�7�Sdo#���c�MJ7Z`v�T���z����C��ϗ�L[8�+��ȼLw��P{�^\�)��c~1"wC�^��G��g�=��IHϣ|��&x �{�igLϬ�Ov�j��B���Ɏ���)1��F�_��<���,������S:���0H�X-V����һK�eרβ=�!����a4�q��27��?�r:��yA�Q��0z��o2�����𾯵��C]{K����3�ʟ��
n��g��ç��?2�Ii�s��l�#�eKe�Zk�_�劽�M2�\]J�1�I��o�(��4��g,�;�߼���$��.�턨��Y�Od�Q�wm��0Ȏ߂�S�2�L�� �w�g�Š��u�,J\���ѻl�]�$���:�<���'�=�|/gi6ƴ�P��n:��^��������M~��HsV>�~�+�J�K�^�Sv���[�D�y�H�]��"�*'�ҵ�J(����`?�W�Z��e ����r�Q�~U���q�n��|M���r��X�X��=��t�|�X4�3��b�&{%A�>�V�h;�nP54f78/�"�F Ê{mЬH���v<3#��Is�6���z����ќ'�1L?�a�$CקFh�;%[�cȳ����a|��ꛬV�p�� �[���Å���|C�쥎�������:�vˑ�����������6�c�lcQ�l}Ep�⓿a/o��LO��i���
����J��KOZh��]=�r���`=���w���Uɠ~���S��C�:��W��u,�X�N"'�u)N���u8޼� ��WMV;�E�?���G�5�+a���Y�4#�|��zW�!�xl���o��6�M1&]�㳏�S���zw-��? ����/?N���
��$�HC�$��1b*U!��)D�  (d��4Ig���{�t�^=�bL($J��w���r��L��и���T�_!)��Ê��Xp`���h>ݡk�?����2;�e���u����pY}�xY�]��@�fɣd���S�`oHp�JP�	d.���nfpEc�3����EI�(������8�)�[�����Z����:����恦�{����ϵ]�H.z�puH(h�@B���"�D=�~������ӯr�Pqm����I��C<�rFj�;�~o�#�|mF_];V�sR�i��픳?�3���cc$NIz�����M���\������Mj������3C&3s͹��v,��jd�Jj����L��5>�5��=u��^?/1�rR�\l���[�4|>�
2j��̓{=�}��!W� 	X<�>J_�e�Ηs����>h����7詻^A�������M�<�~�>��Y�WX�jڠ#xr�צ�q�g�(V�IE,�'�d�D�� �3^(_,ޯ
������c�og��!c�Ċ��b=��0?齗�+SF�YZ�L}��������K-\�o��"�n�c�MYtN��+�D�g�ZM�����F��uŸK�3�� �Y�N>!=���6���0��� G�<_K�ʯ7,v�ߞ��ܞ���oFzn�l���Ls�9�`H	�d����-�����N�ſ���l�� lq|�^hӶ5B�
ˏ�?7k���e�O�b��i?��S�\�\9}X��3؍��Dl^� ax���yj��	=鼱Ӣ��\U������vO�6���6��ѫU}+6�Hү4!^c��� ��'�'F'�\q����\�uO��M���%6����#&�V_~K/g���d^�^�H�u���״�;1^��;O��=�E����M0�����þ\�B����V�=��T:!������qM|'zTD"+��HиAS�|t��ͨw�6xN?�[�+�'�ߞ�f����B8�'���O.�]�(�_Ѿ�E����z�ʼ�����/�o�PD�L{��?A���YEeAfH���GDޚK�%�p��bgF���ɴ��3$7��o�EV>����m<������
��� ��i8}`��|2D��ip>!�Y"s�+cbFG���a_��?4��.�<��>�7����d���g�|����W�4%I����Y��pA�Ⱥ���#7F^7f^����h�[���}փ/���3�?]0�r���szu39����k���|,���U��A޷��L���m��5��2	��W��݉R4�k@�/+H%2�[��ۀ@?�zT��]X3�E������T5�LH�"���} �� �G��!�f��b�US��&�v��G~jeK4�4'}��h�
�h0?�f�+�sMA���&���qF�Ʒ���D>��j��;�� 0�R��δ4��%��XY�,T�% �~ɇ��#Q+��h�E�����>N�|�1��8,	6�6Y&�5\��.�K�Zr�mQ�0��{W�p�EFZ\Q��3�i�:$|@��/�(����V��2�6�㦥*_9|��DgH��R�c���6�m2�;��?7��lFj��3}P1�W-)Z����f�<�Z�3�-���r����y~]�
+�N��H�/~�������\�����������������vS}�lͲ���ŶXm��^LP�G�n��$V_�]��'���l����3z��H�*i�:�k�g��>�`	HgXH��}�PF�z[j��kE�Ũ|��ސ�
�*ԓ�o��7��e	�j����_]h���N@��,�-m��h���Rڹ���!J(S�cVp�ʧkw����C�ٻ��R������#EZ=�B7oc��G�&	H1���ϨΌLɿ��E�#J&� |�qyMTO��J螽�.Ҕ/裱z"^	G��x�C~����Ƈê�H ���?�yD�OΟ���^V�R20��0���_�N��^��y��X�x��>�<��Jcv9w���d���V���Ճ�LV��{�����ѾiAi��8�xy��P'�
j���wF���YYv���,����s��y�-�/]"�.M,�Ç�'׿4�U���pX����UrM7��yG�u��o���E�oH~���J`�y)�����0?I&��m�.��Dr;�q�l���F� �����I���;����MX�[�P!�niaDdm�"��@diuNڂY�	�2��15���O���a�p��%��]?K�t�O�:�	A0�\�U~��n5j��7Lq���1@�&��Q�J��W �v��I�H�.4�찴d4�W�E���C���	_Nq�	ubQ��{�f%V���O9���Ap�Վ��Ym!�s���w+(0z~S��U�bxc ��dl��F)�ה� �o���������P'5mL'-�N����*m)���H�����/k��m��cm�L��� ���5���$�	���"����,c�z������ZՃ��7�k����/&��D�>)ڪ��'.���� G���&ك�Y�zFlT��d����b��^���ue� Q�����hlٛ
�~0a���l�׾Ď��	��ާ2� I�|��"G�{�[_�<������M@!ؿ��,����y��:p�$ �#�Ai����@d��.l��G�2�9�4s�S���=��.�^����8��Y|�YV8t#���ݱ�I���n����/Gm�
��sr�L�4,W��Ѭa�$y�ylP�䪉ִW����a�vЙ_�SR2���\C�����ʣ+}�����J��
��6�+�����֊���"��,��Q���ay#��c?��S��e����z�<����Ut�=����Z�lM)z��nDlY|�����A�b���CC����z����o3_�ˊ����i���d����CAc�<B�PZ" ��,N��������-��u���/��Є��k��n��*�U�=��/a��44�\�ܓ��#�DX2B�{O7�K�T~�j}U&�x5��Mf�7�J����1޼�q`�<H�G�t��K��F;����C ��ƌ��E���DH�A!yi�3����2,��aˉ������yhw���I�8:�q'��u��"����#��K��u��=�>c���_C��`�Tht��W奡70��jF�Z�#�?S;@�)Ы�	�0YB!��Q���I��s��}�'�?sF��Y.G�|�כDV����L2�n����?������n��4��e��]oG&�QC�����<ۊ�[V��B86��le�MZ8�|r�sN�<�ү��I�xW��� ٿ�ge�r�+Q)俥����ւYE�.#AD���P��x��uT]�E�9 j�w8s�;�:�w+�[`4� �m�����:?�S"0p�w�d������D,d��or�DSǇ�}v͸��ƞ5����Hΐ���?+A�L�B����n9"�q�����~�)Ȁ�xXW�<���0gQ�ȘyR�oZ�ا��ȃ��t�0���[J��f8sT��+��Pɳi*�݋X\�Z����س3�v�U���I.��!�Bc�g�H�	P���7go�\^E�挰m]e�K[�[֏!��w=~�Z���N�����	ئ��	X�����}����YG�2�	��0)���?�H:�X���G�Z��R~��mc��*,��^�e�}����Bsx������XN �2�����t�1�y�uÓ�xR��D��{�8W{"� \bI� �OF:qR��`c#V̥S	<����O��og�F�Q�~e�^�wײ�q� �l�n������:U��µ��{�҂u�t3}�)ͪ���� �z��H/'��d6��sH�Wuc%5����m����r�O��Ѧ(6U����uNw{��߂8A�^/�������U��8�{�@�@�6y"%jO83�w�˭��!$s�o�ȏe�Ph%>>V����>�$��:����}�hJb�����ϔ��0�_OiD�ki7�w��f_I}�����r���z���"�c�0O�e�a���u�£�c�ۆ�I��AN��8���u�:n����g��gpuZ���V���#�9�{��4ٖ����MA���͙���\t6j?�Ed ��o��~n0��0e;e�C7�ѫ�3�bG��|�;��m�����!���HP�и2�N�6�M}߳Pֳ�6���|�64u\$�b�DB�v\�$=�*�����q�57Q)��bƈ��"��l9��jsA�(5�����Ĕ�&;oXU���G5����'���]��@��Y���'�M���� �G�0%�f1��pV
��#E� �o��-#��A
���3��H{*E���!�}��Պe�}��w��}�� >Au&�ze��2z�X�T͙�x��m*,}�e9�RM��6}��K}����6K�}����m��wy��:v��l{�-?���/2����� nL�seỽe5L�O�D{pE䯩l�p��L:[:(o�����nM�����(柳:#{��&H�m�����5� I!H�g�ѽ��(�Z��}0�B�7��\m���F��;N��e��u<�9B\��:��%�1��C7gЗ�.�^YaɬQ�\���9{C9���pD"G:����&e!X;~R�<2˹�;1A��\N�~�4����B����MS�]�*�>/x�(�kx�}/i�}5������p�����]KhEĴ��m��L����-����6�1_�?S�r���S����Z�
2�o�M��@��qW�ú��(Q��8&�9۰���v��]���w���.�mR~O;"���M�]�wױ��3)ޚ�KSF����4���1~�������J^S�N�������gy�b?���L� ����L�2Ok1�n�J)O�����cE���"I�rԶ�������,����G?��ٗ�#��"�w\����Ŋ�S*&�[����8�e�����5,i���WÞH3h�ꂆ#l�	���!����M�X�|+R�y�o�~��@%�ގ�!�@e��l<�C��'��Hp���--���\�cHR���ؗ���+8i̘�~;6z���Do��3:���f*8F-�����4�v�ަ�L��|x_���y.��뽚=qu������0���Y�	ێ�k߆��� �έ�	|�}�S�}U�[1��،}	Y���g7��X��柇�����]8+>y(/��勿��P�v�ظy!^��ܴ]�|l��O,��ۡz��O�_��#Ȏ��[$z�ȇő[$b1�����]���^�-�2���0�Seo�<0��F@�!����n���qn�U_�Ԧ�6�Sk�=wszQj ˌR-���ˏO:ĔX�g���= ��@$��Y&J,�Q��5�d�� �J�J��f���A�N��7*�q�+n����9��ߨ��nYY�)]�?�O��$Z�<����6�*" ��Z���H������lz�d����J�wě�~��akϦI�����y�$�̣^��e&�]&����K�s��LEM'��*6f=�qI��&�E_]�л���t2QK��?l�(���џ<�UoT/�+�����ԕ}�D�Ev��w�T�3'�$D���Y�T���˾�C�% ��� h�YT:9��[>�4�(��Ue��ʥ��~bsM�Tı�Y�.G��s�F}����a�B�������p+"�8�	>Vc�t� j����ν�(��g�\�%���HI������F [!���=���(�[=θF	X��d������!+i��_��j��Җ��0w�W��Ugp�Kc^d����
�h��駴d��H�O=4=}�3�\���za_���?��]���Ec�ڷ����a�|ww����q��b)Q�s�7�����;&��%�'�z^�J9�2'  ��X���뢱����?��4?%�����+K�jt�|ҷ�¢����)3�l�`�#��nQ;dKM���`�F/�3k���*k�`�,�hj�*ח�3_�#�I�����UwӔ��ڲ��`�g7�,U9���}��>a�6zK��w�Y7<;|\&�7�ʶ��)��-K$b��JToA�����Tٛ����Ys���̈B��=���~ {���^YCjX� ���Z��"���`V�i�q8Lک&��qn��T�[T� �>qP�-z�>妊r<��G6��6�7{�M���y~2p6P#��D ��<��_�f��nE`/M�7�B�����Uz��|)��5�ԙ���2Bu�qjN[�F��iN���W�x����ߵ�_{�-9a��n@^1$�4&]�PM����/������C�Z�����+�F� ��o�'����D/8���l��0J����`~�ӛ/���N�����U�QV�O�~����Vvl�������R!�O���5�m������!18+Sm���9o2�f��n�:�:b��e�����Nvс��n�4��l� ��s���	���|v��&�W�!6n�1W��Os0Ŋ�d���3O1�& gۘ�W<Q�P������i!(�HNıQ�ZFըX$a�#��.-ʇNH����K�
�Ԍ$���~�W�0���9=@7��x&��Q�T�>Jgk(L^�mM��;�DD}yԽbjd�=gr(�:_��&n�b�P�,㤥����T����'�P`}*�q0�<8�?�c���IV���?���:�~�/
8U/L`P�P�,s�M�z��
ȟF�.&3�����6'���)�19��2�9O��B���/? q@˸�z���+2�1�z�̗�l��wm�Ң�P���q�03
�k#��D��O]��p�Q�xI����)n�C�Ήh*��ȥ��J�}UM�;C�Y�{+��!bza-���0��h�*�kGS��79,Ä�b��y��j�X���ω�3n��j@�b��zL�G�?4ƒiK���C���-`��꼱��D���NV�w�a�[��� ��=V����D��%Z��*�ٚo�o������X1{p���K>�w�Z��=$VXt���/������#;(\�]��|Z{��<�&b�um1�`)�SD�`s�Y�K7y�SX��EtxHpÎf��w���Fn�\]�̾�h�9#F���u��)�K)	ʫ�����\=�J#8� )~���r�C��O	D���G4��:�Ÿ��2/�����N� �Y��Yq]���0���
�&%ڎ �!`둴�0'�nzp�����*�2��𣇅��齼[Q���jCX�L-�C�猞�j(Q��j@�I�4��;��Co�C�8������4G��&#H�U����gC��*<��ǚ�����T��^���V9��l� �`:�|�ې]�]�ݏ�X)�Y��h��m�UQ�fp�)���J{Jڳ������A ]�E]Tޝ���v&+`�F�oXԊ\�_�c�o_� �X�������-�O�
�|oq�}C�kɽ6=*�l����I�n�}����t�2���_vx4�T',I6�|d���y�$��9�3�F�wL��$!�O������G�~KPÓ`FO6�_1�/����)�x_�P*{�B:�3i��r�H�&��%ʂaM�q}�(ˏ���������8�\[���`~0H����l��zm�h�>�3c��/���3~�K�C��m��-Y5{��������8�!`��|�6�{hͲ�p��W�eβ�n޻�/�o��J�j�=�n�p�;1��c���~�	��o�7N�ʀ��A��~�8S���F�$oK���ϣXb��9�[ף�/�}�����穋U?Ǽ�Z:g[��!�W'�҈t��b=��E��Gg���B�afB�K����N8�����K�6�_��ʟj�?�����j/y���o�Y�r��2�%�t�'%$ju������e!cTjV�����[��0��#⼔�Q��ku��bJӯ<�}�_5n6%(H�U����S��kpU�T��Z�J[�J*Tx�
I����B5�>l2c�K�qt���@I3~L�)=���Flm"����)6qW����DB '���+�E0�U�����63�g~7�q,��)������,w9k=A�+�X3�ճ���H�C	Q jZ�����Xa`fNxy�8�w����x���bdk��~��i�&~\��ћ��*�Y��g�4ڏ�s��#��g9p�T�&�t|����%yI�ܔuI ��ߜ��a��/j#�d��R&Z���f�V���N�!�xR���ef�N"Vƫr�!��A�}��*d�����}~�㩏s�٠W���~�����B�u�C7@�m�3O ��L�L#�`�FJ`}\��A���2��� ���zv4C"�}��mq�C|�	��2\��_�EK��rZ����`��� ��jAR>(0�H�dL{�/b?�o��F��ٳ�-��w���x�`���K�����_º���:��V+�F�XF;��i�����Q�E�p��������D�ߦE��8�
c�M�C���w�[�>
%	l����ڜN1?o��l�ڗRe�WR��^������9�_*�s��ޱ��z�G:�X��
��_��˚��|�d��Yx�>+��+jh�-J�ӚJ�agҤ�#������v�}+_{�Ï�����#�٫�����A_#�1�2�Ai!�$�+��9[�Rx�d���^�T#CC���;��nUt��2�����Z�G�0P��ʙx�Ąf6�1#,��B2�n(�f�i��lc�����	��~���l���&;h�*�`��,9�
�������v�!!bJ�  ��.#sRL	�l�g�\��O������(�^�&�`U���57Q��fz���4͡���z1���sFe&�Ⱥk��Z[�ݪ	8d���! EO������j�:aǬ��v�y]~�}p��5m)ۍ��J�k4f�(I����n�֑��պ�i>�I�?�r4v��X�f�œS)>��}��P�
���қ�4����t1���G�[|�_x���[ܽ(r0���`�|n�C����ˏ�����L��._v����G�!�V�(I\� �`X9�iZ��ሄ���n��F�r� >0�+�\'Gz#�C�<�n�[~k�{��SR������SMY����wo0Ak0�`Q@�,�Y�T�I����o�]7�*n��v7��`a-���w/�b���o|�_����k��
�87�S�8Qɘ����5=���'=�;�/�T#�Y��#��S/��RB 4,��ۑ��-�8��b����%

����hn��H�ΐ��斴Mѱ�5?u��q��TѮۍ��3�쁩��]�ğC���ݺ�3���&�L��P-�o�'$�67��6��j��gΎ>��9?wWy�OU~�婋K�?5<FAd+���.컭����������T��SS��𩫯����ro��1:�XD-�]�=���8b�(���I�����<U6�� 2ig}����c��f;�z7��w��A�=X�̛�m1�}��E�Cm���5��v�2W?�F;Ţ�xz�Q��긵������nX�،8/�F���(-��`���"M��5��>�q4��\@AB*ߗo�\�_��Ew���6��]�k�'�:D=��C�%�A7�`��`|O���7�H>ӽ�="I�Jy�!*�?!�����c���~, 76vU8p��5�I ���w���Ȅa������4�Oq2�}�Iq�J�%H��y��P��~�����eG0�g=��p c��˫�f���ӧyd�p����Ɣ(���v08�5�������Do��S�a��tM��ǹA��o+���o�2CC���5._���m����~��OI~�[�^�>��i��czE�'�	$$���oۙ���c�4��=�^�i,Tv�H'�S��?)I���ԜyƘ��g��ps&�k	�Y�c���	��t*��n�ɓ�PS��$t6�~���liF{a�㝽���G��Y�b� ͪK�Y�o ���ak��I��S��m�-�L�+����P,���_<Je��=:}���0C�e%��ٮ��1�y��m� �	a~KBSJ�gZ�h�Q㟹��#
�\1���,�� �[�>��WQ��,��������UC�<ܐ8kL��(m$���ۆ�@����+��NB�c��pKX� 7D�ͧ%!F�./kl�>���m�=/�X���+|�ԔL�)��g��+ׯ���c�o��*ic�9h���2����}_=ж�ǂ���@G�X�
�S��9[�i[��޲j0%�mR˚����@)�KV@�h�������G�WGE��_�0t7HwI� �!��)��9� �� -)-��1��t�tH~ý��~k͚�gN<����w������=v8!J���P��,���u��Kv��˔4eR;~Ϥ8�:d�=���+�U�h��<�D 1���V ���Rl��S��7+aD��x�u�NC�h�g��{m��q� l�c3�)�C[ep��H�?E��Y=�k�S/EP��l�A1d!�k���=j�8�n�	Ω`�IAe�W��^��.$161�G���:ëw��w�HIc*�e����l�~��a�YwԸ_���� w���3��(���ё$�des���P
g2 �,�v	��R�3�6�^!LBC�d��n`aЂ��0f房6Tx��@���glJ<P^I!�Jyd�4%E�uD�|\�p|��ln�p�"f��g���e�fJ�b��h�6�냮�f����9����K�7���e �K�d_���@~��	�6,Ncܬ&\�J���P�+���V��pRt�8�������e<������ֱk��B#��.%%G� E5���삹�wP��N�FX c�`N����_!�̴�Z��d+�ɵ��O�/j͵e��78I���_;���� �gW��s�����wܬ [���6"hH@W"�&��LT2-��
��RB'i��.R�'=�,��+ j�u�����ii,U��$��N�������jk�P�q������N������c����|mqb�c~����63]Nr���(� �U6��c�!2{j��aZ�!a��%�U��pY���޸���0%��*eE5��1vJ"��)Ղ���2ָ�J�#������ͼ���~�[�+Ų�1(��`�2e��m�pS�d�5���^E�}�E:�|if�)Eu>}
 ��\�}[n�Zܥ�|z8j�h�N>���� ����E[����h҄1�J*�
Q����}k�o�b ���%9�z�	���.:�a ��IO�s��H������&K������i�/Q�R-Q�{Gi�3^5��Q��cR��~�����^d�m~����N�#�?M3����'�g	�㻒|�u 1|?�6��d���x��N�v���e>��N�wR
M]4.���{.6����4׶����5}�U��� ytd���My4���j{ ��'o��֘q����T
�`��H���%I��9�;��7���q-W0��;~|G^�s9�s���sv�����؇��r��­�̄�t��޴۳!��[�U��b�y�"+&����k8y9�L7��r9�B�Vk����6����iC�m(�����7�^GQn��@�+kF(3!��J�����XV�����Տ#>�x�\�*������y�?�.�D��r�@�@0�"J#����*Ս8.�b�ig%`��L+�py����ϋ7���Z��c���<�yV1 �����8�8E�oX����@bRe�F���-m�}��GF�S��ʉ(��-�b�#����P_3@��9j���>�j?3T	@|�Q6I�@�K�gF"��}4+�d���qᢋ�\o��|{&G���@�(q� c��D��%j ������9)w7D��ŒD7�فut�}�f{���I��'��m�T�A�FF$
�(�J�O���)a�J���;��Ǧ�z��Ǖ��=��Y���u��n�ΆFΆzZ`|D�[*__��in��-��L��L��3�����'�M�K�q���j��b����ņdA���w4��߾ǲ�ո�� G�	����f��,�W�bߓd��('�G�t@\^G��В��&�f�r�Q���uۊ�X�����9���-��%�h6#�tI��a��2�	���v�
�I��(�9L��|]���>	�cM�z��?%�پ�����d�;c����?rn�ڨ�{zL�F���;(��o�$��̑oq��9N�4���s���9$%qש�Y�B��b���{?��<�7��*���ļU����}�	�G�2�#k��{���k�ǧ��Ѫ̈́/	�X�V�t����x̌��-����%4�(���*�`~j��Ɗ-�z�*�֤��%����V֑�l��p�7z9��7ÿU������{~��h�U��^�~L������b�\l�����C��B�yB=5�E�����K���z���k&���8@�R�G����{&�u�,3�b�n7���e�kI7���	+3	�X/���j0�Uw�j^��ƠH���<���42�\*3� q���]���l/�!�p6Ņ+�[�a&Gm���qӆ��ǲU���ܫ�A������X)���ݙ��	�Ց��z�;�1-��e�K\
����o�p�4 xވ�L!����ܝ�=1�(�B�'#_�!�f�(2YZ��o�_��e�~/u"koŸ��z0��*{<�A�1э��u�|�{Eă�	G,m�H,��=]ȍ����}{�F�@z�{f���y�V� ���^B��v�޶^��(�a6�DC-�/+��_��|Y��8���\ty�yy�á����z��Ax�L ���oE�k�����+_��I�'�56t���ldc�9 J�	���~C���� rPq�F�[��V�����D����� �l�i��߳�����?ˋ��¿��e�oL�b�r�Ո�	�ӄ��0_M���O�o�hͧ9�$Q�=��<Q���i����s����p��Ƕ�0�
\'�oЦ�Z���+�Y=�,oƚ$�魡�;t@VP�-�/+�KA���g)Yb�.�QHg�����c����
g�Km���:Y��9�.�.��53P9x�Zϟ�kr����h��fk4S���R>���a��n���v�w#���vޖJx>_�B�0�=�j8�O(���v(�k	�y�oko2��!��|�b�zz�ɲl=��ߏ~6ե3�����y��[z_%!ü5(����L��9��J�����S�j(srw>���V$�e����������SK�ρ�Y���}#��6�&���ėo�eF��R�����?9��·U����知���7j�ng7�z��7�|)�=>��3a~:�T��K�C$�jB�yo��,~)0��
i���/���&�.�����k`.��w�RG���r5 ���)J�/�]-7D��s��(�l�k����@��J�!"�m�b�JVj\k���N܈J/��M�o#*�OF��7/o�/k�p�1Y��DP}2 �4�j�hw!@Q1�y'aղ}5�&�ؕ��i�z��+���/�kaljG�'Ejbs��Cc����a]��]�I.O��|!����L��q�2�P��|3�C�Ҧ�Ȥ��e�M������h f����X8;�X8۽h9ۍn9��Z��'e��?px��}��h(�wR��@���O�&���M ��Ii�VR�'F*�*ZJW#�N��Z]ue�2$�	��B	F1|�/Я��}3j�ѩ4j^o��M�8[����8�H���̖��E�T�|��w�W<�Ϥ�對7���l�l^�	E*��2�ô��A}V>��ѝ�b��^�B9Ό���[���i�i|���μS��������h%��{p"F�9+�D�X��Z��~T��7!��8Kk[�P���)|�V]����h?��z����ʯ��^�AD
�E�R[,fv�O�p 7^.� �)�pكM�|�{��S�� ַ�}}����w;J���=��-���l�>��x�o�"�iH���+���	����P��g��Цv��
���8��ۇ9�Y�=�Z7��{������<�d��Sz��������Zp�FÑS�x-f�a���Hif��[�:��L)��0�sP	9p?l��X���M�s�L��|�6N���Yb��I&e�L9��P�l���o՞��$<w��>ߔݮ�m��m�"��GD{�2U`B�R
З7 Ɔ� ��C�\���~��"h�d��&A���t��O����@��� :�`Gftg��-���(�?>5�\��UP6x�ce�uG�t{�(лEK[#_�ʩ�z�%�C[A ��F�퓻@7ejAz9�:�`���@��r�&Pca���Cb`dN��Z�d6���o��Kmޣ$��P8�opZ�'����X����tg�<֬���-�邋�J}�J�����]/�d��7`��y���������d��̙�Z#��Gύw�̞�O���Y|�_+����ճs��%.�AW>�x������G1�>o�(���y�5X����٦�nqZz��������`��#0�ݖ� �7(Hrz�,�������~U�� ���#�G�IskI�Q���t�!���[�H�Tg�-�0U1=�$�#J�r�)�}��yY�	$Xg,C dG�$�O4�j�v���k'r���_�f#��#͹�r3����⦐�(���o��k�G&^����ҥ9�B��"�ƛ�\D^t�Vtj%�*)K��F6E���{:/����\I��(w=��;_��Z���[�j7�?')����t���bO|�5�Qٞ �7��[�����DKa��"埙S�����ӔG�2�X�M���i�ߒ$~�R��/��-����,#A4�,(Yt��7'�ek����&2$g����K-iG�#�~�l�R	(6���U����Y+�a��/[�,c��:1#��EОoA��.G�jH�@��#���)����2���	g=���OpJv�G����-!B{Z���h�U4"��!+Ϛ'0Aǡ�f�?x$	�vL��6E�?���Mw
�!�s��w����i6�yz$�Ut�E�J�<���^B!�'��ad,��('����%�!���Hs�Ui�n6r��r)w����e��N��~�~z.�;��g��Ū�d�7'k��O�綡��K�9�Lj,��>	�>
%�:яc�f0�����
U�x�?�4�P���c0=e�l��`�(�x�b�XL��4���9�3���N��l.�c�V�Cp5�=pkl3��Z���y���[��X
WZ�����i��E�@���$��%�^T6���G���C������^�X
n�E�e����,3/�\�?��.̖���f7�è)_.�X?������Z���!���F�zU��oP��^'�UHf��ňi��L���Gև���&��+Jb{���F�}�}�D"��r�q�#��F@У&uc3��2�d�tؿ�4�8� �L�������x9I?��q�t���Zo6D#�섒��p��cQ`�V���a�6m�oBG���!�f@�G�S������IJ�|,��|�����,�V�9����k����V�M�ٴ�Z3✆�7��S?Ƨ�r*��2�n�x�l`����>I3�-	�`d^����@(2���F�9�%L0e��#��YI,��&�z�lL����&B2�0�0EʉlCkX1n�5�N�H[ڐ�/d�K!�Մ_�D��*rX�V�*�:4�B�3�,�x����߉0�n���2A3�l�>d=�����%p�E[��
q��5�u���n!��l�TٝA�Ϟ�34n��������C�j�X�����>~Ѩh��?Ǵ`K���O�G�W�� ��(�~팿�DX������Jwza����I�ⵉN".I(wݙxU�������6Eܗ��ב�s�qw��$@ٸC�&\64.��
�Z��]v�a�i��S!_�n=��E"�e@*a��Sa`��*�=��m{}5�J�%�$�������d���E�q���rC8p�D��V�
-��.�\��[�{ҋ1>�k`~�	H|�}�Ӄ����-��n�"WuB1�EdF���:%׭��B���I6���n��] �I��8���%�I�����t��q��m|6q�i�I����#9%�Lۼ�ٞ~Ĭ��"�S��4��	"&ptbE�ߌ<~cH}����\�Q���#�[�h���A��b��tD�Cn>�G��U'j��������"Wn{'��9��՞��|T�Ò!SN#uڳ���m���+�Z��S7Y_b<�y���#x�$�-DA�UI�1�*��G�g��LH��� ����׭����:����[pN
��ի��֛�FW��4�wr<$�]��f�aB�f�ס/M�Z�T)��������N~�u|UK�P8x�3��
�����K�	u�=���Ss�9�ƲSPH��U"��*��"qu�ÛD��.��P>���tD�7��&��v9���A²PV
�tz�7��9~�����d��cL��@>#+?%D�� U��'�h|�C���(W$N��؏G[�2��+l�vtA��$��(�U�=��v���qr]'���E}FpZ�,�>�HW�/q'-n�WSy�O�u���+��ͮ;�&-n{�Z�Y��@NuadE�K�&MK>��	,3sj^ a����t����T���TPl,P��6睲06�Mw�4Q�N�E�+��S$������,h���I���1����4vƍ1�I�k��&S��gi���:��b����p
[�O�aWR'���GE���u�|1'���D�����-��>X=hz
z76���u�2�!JV-�ҟy6�\�k�{��>U�P9��������w�lf\���(��@� 	�.gh��l�;�hԦu��zǝj�O��b������V7�r�k"iN�ױ
�\z���O}���0/��:���^�pt9/;n#��
��Z�B�Z��2;�|]�-X��l�j/WY&ʂ�����_��Z����c4��Me!�sƸ7��[U��|�v�4�],�G��fK�K�Z��DPyaD���C{8!���)���XI�f�]��*w��Y�J��A��2���n�_�	9 �֯�I�G�!�Alr���
�D���m�H?�`��VOzB0��Q�/���=\���h���	�����5�r��i��1�dX�	��X4�hR[P�X���K���1<����Z�M�o����k6�i�3��:RV|C����hkX ��E��">EN[8f40P�IڅR��� m��N�t�I�ַݱZ� 1im��,?~Q��i6W�'ʟ���UGT����5W����?jXAC����z�e�#?�t�$��Tu
3L��]�ӳØ�đ�����*�&��>t;�w���E�V�B��OV\���pm= ()�D���aha�?~�O��5�j��h�;"m|%��V=�d�a&~S-�t��np�;�6�啸���M0�5
}CU8��-V�dO�jԂw�i68��h�� `}���%Q�V�7�W#,m���-Nx9����7��_{�!��r��b]Dx��^�m���Q�N�7m�64�%% �`L\��^����6�O��|�|�`��~�Fڰ�]9��#���pez������s<Wc9�5�j{����b�I��q�ᖙM`:a&1�y7W��M�V
�#W�5�+E<(I֏P-��s���������	���Ӓ ���or57�4�X��[$��4�3����-���ؙ�9x�nҼ�?�2Jly�۠��U�H`퐡�/�i(Z�D�C^�#G��VGD�
~R�`(��h>H��Gފ�K�7g&��}�f�&Ĵ�K�@�s��ܟ�su��=���@<ƪF5J��\�l�@�y���_/}w�����l����	8B�Y���A<��c9�+�>6L�.��l'��w����������?�[{n�8��.���Ɍ����t	���+�P��6��Ԁ��U��6�--��wQ�Ź�¥�h��	[]�Q��!��݂��:a��:��Fİ6�^��U�� n��փ��@������'Z�x��p��0�j܆�N]̟����m6��7b���"�2�TG�o7�ԲH=���6>
>h̜,~��h�q������0[I!�}F��a{��=�M1��oI@��j@���7sVA���M�&_�&y��̀̍�+������30�~b�e;͞���͠.E݄�s���-�画�(�Yc}��⻜L^���N��Uxp���K%�,��=�EUPj(|'��|� W�L7/oLZY	�U����W� ��!���@`3�f�����t��\9&�zy����W��}	ṕ{�:�tO��x�|ٺ�ZS;,]��w��激W��9����)�� ��%��<� ίsR1C�C�0�o�l���@㨭��[uk�ͻ(m#y���5#R`wV	�5��Gs�=ɕ�-�#��ɝN���ފL�#�����pL"�v��'����`zwJu�j(���8��.QҒ��Ԩi�ҍ8j@�.���Plr�Y<����a�������W�]�~��æc���0����;[턉��^�Iq#Hϱ&T��˞���O���$/!���p�)���c�cl�9�қF�j�|�<$e(J{�`o 1/*�ۭ@�M�& ��e�	HBE�"$Qt��H���F ����i�W��"�7�=3G��S��:�NE���nz�~w��@���t׃�E�f	vt\H'Q�1 ~�j�`#�Oׇ�C,����l&?����I���w�����7���GkV\�����C���S]A�0�Z�ô�H.���i��I1���	���<{�ƕG�Tn0b�1?����YI���\#�;áH�9�{D3"ZX���uS��-.X{W&��C2�ч�����v�Y�տ����j	C�4��l�xq�՗	�M�诓_��Bt�4)D��Sl�cI�$̤卌�мGPđ�"�c��3�ȶB%�7cMւ?����9c0n�0�������XB ���2b{$vڟ��d����}E��a�F1 �R�ą6;�e�x�^�&��UX�	5�_��K�k� ���<��� Az����)k��!��a�K]��f��h���|�&D]N��^�9<�T���{w�+��R���R������/G�}LD�V��"T��a�<�M���륹�-����^{~`j���P;������8�i���������, X�B�1c|���%C�Ó�57���Æ���PX�F��E��F�]]|����4��:O��Ĕ)���d�n��S(��װ�,��o-	��n���O06{L/V����}� ���#��=�1)3��m�o3�ۜ����z]MkP�y���m�m4v�j��{*�	��:r�o���s�U��B�x��y�l��rs���r��iı�G)d%����5ԅ��ޏ�Z��K��:�JN�UN��O��)M�#�j�)K�9�1�n�T��v�L�VC���޴��'�'�6�����K����J����Y&-S��Z����(~w��}�1K���|D���h�l�'1���BH�����\x�qd��A͇�.�)�!�p<����1uqŢ�V�\^u�̊��ȜF�Q��S��ӈ)X�Q�@f��tN�=A��[��Sc/���o5��6�7���f���;4����.�:Fq&,FH횧>�ƾD
�����$iب�������ʝ��B�B&C&�)����-`�?�Ex��4�<�MI�_�,fk���L���aEQ ��.���u���^�=�bO	҇Kca����y�9Q^긄Y�qS�B�5�
����%`Ru��P�A���ӽ��0ܓ	ϡa
��ʐ��D�������HV�?�_�B-(��;�]$!�B>!��Η������6�����Jx7�Wǘ�y;�"���²�� >���3i����۷
+f�L�zdC��;�w=ipw��-|�zM����+��7!���N,�-�� �_޲�����D^���,��A䜘y��B %�a��v�	#f.@�	^VJ!=�.Z�j��d�Go8r�&�'��y�9�a�2��zȊ�g/]���;K"�Wų5�D���ȫBb�
nӥ�jg�����m�֮qr^��Pù���}|51�߱cPIji�F*�Y%�  �Ae��]�vI��S�
���u���>�B�
����8kA2��C�����{����yBN�WT��T�.E���!�.��mE��[�C�I��K��M�ƪә6H�Ч���*h\(�İ�<�����}B���}��ʮ+�IԘ �a��匞�{8>�[rN�����v��Tj��Uu��J���A��{:y�,�l`K��|j]_!�_��]\�{����|������{��9q/I��+��(7�v>�Yb�}ɬpUj�{~;�"L�8��bd|%�r��|�S�:/���o���.#���|±��[yG^��ѣ ������ *���%hߛxL��O~����
j�>���VW��acA	RC z�����>4�~v-"U.�jt����E���	��I_�� �Y���~�$�:JY��U����l�~${�\�7�I�߼�1�ߥ����gx,r�3���A@@�J֚�M�P�s7$�T*4�V�lL�anD��	�:=�w���?%�)�*���NT��T�gPr���>�C~���_g�/����V#'���i	B��ޖ�oI���k��ѱ�lM�`��*�q��+�K܋�>a�%,����+�%+_`LT1��  �����ݪ�yE��
�V�,t�e��kV�L(�
�n�]�����"��;����s�gT���\bc��5�K�c�Z"�v���0G3 {��~��R�"�r���IG��aٿSձT��ƨ��!������IG?�N�~{������%�f�K4�Ba��s�S�i�ҭ��1�޲q��3BCV��"a�7��*��^P�G����3��'2ka���cעIy�?"q0V"q �K21�_���e��˙�x*l�b)-TK��U�����;AN�-؜�����4�{�R�Z1K�L] �A+FdL���݊+�����B�);A��؜K��X�A�T��!��f�$oe�D��6O'Z��q:�֝�� �v��=r��N6d���(m�������h^�3^d^E�>����ُ����a:\t�lx6ɞ4�#�����2X��0�Ib�}Y�&|����e^M'��6�|�K.���C������&k��cG ���ʠ@6���0�~E���9��ɭlﹶ�Q��z���{�v휜�[h��H��=Ð."�G�G���qlX��w����+`�����u6�I�\��	6�*�ͪl{�mT���Ĉ,�n_�!��R-���=zS �E��B)�w�QȽf��d�QQ�^IH�ڣi����Ѥ�1u�1�_�P1���5�O�~̹ �f�i?6dx���F��e���R������\���X���������w�1�� 4��h��Q�ݧN��c\)���naa�9�Q���wY^¤ȟzǛ���Ib{�����MK����)AT]�b-�F���byn��R�j����b��sq�vA���psiL��R���#��/w���p(mZ��|G��@b�Ѥܔ������	�>MV�ϵ�_=B�wA0��^�.A���s�ՄI��_Q��C��lI�79�X	Jo���o��bMJ��b?8c�a�s�QC����ޓ�B���v5�)�Vf��^-Đds[TE�=�_o�>��кl֧u�V�+�\چ�����5$�W���Sݝuئ��#7H��U���o�O/����D��c-�����]����cy������~Z��bry�z����H���͘E�
k/�-~��'����5�)�f�R�$�0~Y5c�ƿl���".��o�bg��e@9��.�-�%
��b�q�171Q�/Z[%?잪�(��a��˿^�"�O>��Hf5�M֡�XW�/�!N��Ŵ�*����^p5y47�r)�7�����^�<%�3'���P���<�"����3?�`ʸyT��� �1}ܬ<	�P5��f&��R���(X�a23"�Fgc3����Jx�j�I���$kG�s)Z<��v�R�P����
� ��P^�T7����r�~�|ʑ}�FkZko�%��v�:r*;�j��
	oR���˶���� ��G�����:^���6���;��Ǎ���{Վ��"�5�ޓM��_3e��B+����W��:�:gVXY�n��H�q�ͤ�7�J����֛����e����w_.7Og��gɆ6����(/75��t9uSﾔ��,�&�sD)���+��7��8N8+Rп��*)0j#���'<��'\�W
��L����䲸����>�M�TY�1N� :��#/e)P�d����ē�$'1������K�vj?aS�¶8T�����3x�d����Of���R7��y�z|s����!rb>�L }f9����D��q�m�����p YU�
+�1�&$�s��ye�R�FFo��f0.ПN/�r~�II9�+C�Ѝf&V�ޝ�[�Gw��d��+[#G�B�����m{���[@V��&t��p�i�����M����9��>�_&4�<�i7���w^�QM����{[�u��l7�1��C/~ĉ���P����{�e�����k;Q�	� V��U<��V�U�K���1>yn&��ǢI������j=������T��z��r��[�T�������7��h�C��$LI$bMz���Oi�E?NBa�Z`�1�.j����k����,oir69�a�J4ÉZ�;^�FJ������$,}�A ِ���I��=���=�+7����t{��Jp�A�L�ԛ)-R.���f�<�g�*�<�>�k��	�Cھ�i�L��g�KZ�ć4k��%�C�kRʐYpA坓8�Xx4��X�ؕ���'Eq�<�2ei��6* �CI_�&
�;������j��mȑi�W۱���F	.� ���%^��us�~�P��?Q��������"��'0�S��1ȖMY��P[��)�z�F$NT�	����¿}׻��ɺѽџ�0�G������t���w]�Jk�~+n��6��y}'�X5���x;���"��ݐY:+�Nc�֨RK��V���gˏ�i����[H/�@!�"�k,�f��.�i+���3��TsF����!V%ͷ������8����֑��$2����b2�����qE_8 6t�X���F���P���R֔5����)aǢb�#�'�i��q���ȣ������%:!��[���-����ۙ-�� �V�,Nv��)V�ޗAsJl��ah7� ��*�� E<\�S���j�#���|��?�b�"�� $%�L���qz���B�I���� Ӌ���9�Q�b�Ud8I2~)`�����A���F���PX������DUa�`�\�"]���:d�~5�J�����Y?�'��vAp6L{��#r�����Z����y(7�/�_H�n^R����B��ս�G��4���h����7�v�`-m���ʓ#����>�n�>�K���T!�٦=T*\}4�K�{��5�ϼeu�pᄥ��g.�@��Қ|���n�m��;��ۿ(���3�=�8�8`���H=f���$D�a�,!z>���9�0f���'Ո���ʩ2<�N:/[���ܙ�����L�X\Sxt�svb�}+o�A9��{��!̾X5��!2�AI��u4y�i�A���f^��-��˺}�;4x;���L�sPN��*R�!�Y�N��H���"�r��bR~����ŏ��e[�&��\�/�|�x�4nͺx=t�o�~#�+4��ՠ�f�����|�5�&n�E7}0a0/��~c��� *�%-2�/��1�JX\.���N��*-؈w� ��a�Rf�����O�b�����zgV����e�]�F����'?�ܓU�b��t�=���H�;l���-0j�-�%�s��#l`vLg�@V�5�_'�9�DH��"�~�k�����F^�O��!����N�F�T�B��a ��Y�]_�DI�]	��˜f��R2]�[�By�����m?�^�p��
����['-.���3*�P��S� 	���R�K��KE��vʚD#ԞV|�P�L�[e��b����Q�W��#R����c����5Jy`����D���>xCL,��D횿�,5V�,�u����W$s,��LM�<���i�ڵ�E�s-��W6ԛ�}I[Q���$��[��r���I� '{�O;��@vt�%<֍7�~�=��y&�,ޯ=y�8i�c��|�*��v���xh�i��tj��ϱ`�1,8j!R����=+�	 r�r?0�t�T���9ͩ�h��)!?�|���N�+��
áz<���9\ڋ5b�*�"㖈�n���i�F�lrUU�Ú�m
N�xW����(�L�A���'���G���Z��^ �c�r�Fđ��a�qo%�(M�29� ��@`�kǑ㿨�-��سȬ�ٻ�ة�Zn6kB���]�Dh�}
�b�A2ڨl�_�E!f�}dp����p��:�8-��k�7�ӓ(��&$@'��� ��f��@/]wO�b��9/_��7����褲��+ݏ�m�jFl��(nƺoŞQ���iܳ�0��F'ֹ�d�k�Qz��d���Y��rܓ�2yF�r�/����.Y���-��s��b����lQ������I�B���VY)yܺ�2�z;�l���A1��b�����y[9q�]Iɖ:�r��p�V�!��{�m� ��ʍ`��o�Z2��=ɚF��"��P�	�����ѠG�zc���4�0z6b�H��S��'0u��˷"��"�Wexw���^c�qv���Ub��r$���+�Z�c�L�	��4Jj�z�^�	�C��&�e���f�ʘk���Ѧ`".	����l����R6&t��fC~0f��o�D7:x����~|���BO:�F^o0�<�_���Y[��3ie<�c�U��7+Ҡ3f��1������5g�{2��i;��"�;��g��oT��I���~y�W�i4����e�FM�L�.T{�
�/R��Yߤ�u���l��_��'��bq}��NQ`�E�"����n�O	��������,<?���@�l���[Ec�?�0�+_r�۞�3��'���~�n�NQs�(�~�=�ݰ���]���l�� ����+����z#-iJ��2�lq�\���z
]�?�5�?�5�"?OА��^q�_ݯ�Ԭ���/6������'c����:'o��y_O�X�<o���p^�~
��`g�Ý/���P�/��"#_U��+i��B���0q+�-ȩѾ5�"���Uw+���ĬO�5�R%�Ms/|z�<y����:lp]U
]�02/y��Of]G ����_�\����on
�C��βCs|OphX�o��3sI�}>�D�i6�T��#V��}�e��[Xxqʎ�cB���ƮN��ʹ���#��pv���^`c,��t1g��Fw����B�}���7��X! b�w1����З��"���K�.���ѳٓz��ꩇO?���W�97|wL�������L3�9�df@�KIi;�T��DbhՈ����It/9\/�i5��{?�a'��3�}���x�g����ySBw<ƺh�6�e2��lu������B�r����z
���o�,�\�jI#,>k��{��Z��^�?�^��� ���YOj>��@�o/슡�Q��[�d�����q���k�F៻���
�~}ŧ.��X,Z	\l�;�gÌ9g�w� �К:��p�Շc�D�ɈNQ��/2zt�<���\����g%��.'P��&�Z(���e��B�.��P��J��z^�#9�ٗ�X�F��nr��_���ȝ�#d������g��}�`�~&u�,��LU� �������<e�,�cnA'�����֓����E���V
K�E��*g3�+���
��ƒ��3��sfS�\�#��b�bך�b�]�:�ɶ�<�3�l����1�o��ԝ+��z3��B-��;���r-�T[S鍓�&VL0D�n~��C��WG���6�R�k+!�]����%Q���AicK�R���zc=aNGf5���Ga?���YgȐOά�cH����0)c�;�}.;������(r��$�����H�TOK���HͭH�����B��P����"���@�D �R7A��6�fk-��<�kԈNx�W%��+��8]�-��r��2W�11�UW��]�&��D�}!�W�P�0��z]r�"S���w}C�xT%
�x�̷�`l����r�Uq�Jm �N�e����>�z��o���e~�@�Y_�}�$�a����E->�۽@+��t�O�Z�C�E�&�}F'y[���*� ?�E���(��
^R�X#����6WK�_� �Q�a
6�!
��Q���������}�����f�'���N�ȇ3�j+٨�g�S�"����
�["a�ﱼ!:~�6�>�e��e����H���3R��Je|<r�f�\��򯽏X��1��f�b¸دyI��"Kp5�)4أ#��
~x-;������FY�>�Q�N��b~1 �Օ���{,�r��\`�|�|�K*#$NA����b��=�Du~�O�6;��� �� 0��w݌��u�����a5@�z���
3[�w R��wS��7��+⩘����=����߾n�0���$M0w����UD�=�]�Kv)��n�.�rA��.����;������;_v?���9��;�̨/S��2a��N;��z..���C�_!����ǧ�����$�*��qjg� #�t��f�M���1�͞S�%Rl,2C�7&��T�8JU������kt��i�� �$ U�0��s�L+���p�_o�&�
�U��Y� �	jRf�m�Lu�w6̴C����ӱ�_8cM�8c�X�ZT��U�췇hd���6S}���~Ȝ(�}.���':#�,|(3
����h���k�vyDu��c���ݙ˓OC�-���O-Dd�5 �
ss�hvt5�����iV�$T+����|���B�}����R� h�hi�t��l�y�KvM����Bf��G� ֎S��o|���r� ��m����u\�]%�M�GZ�~%��}�af��\��1Հ>D#��WR>����9�'�'��e'	')�Z�.`/;Rat��)�Q�iE���KS�)_3`�dv������ �i�F�w&�G%{�?���K��Y�%��g.>�t�����G��u�h��&LCng�oo?�k�~ٌ��8����m��p��_<f���U_��vd�}�HOq���z���B���;�T�,��3�x\f�o�
~�W�pd�JI�V��ԞisT�媨���L���t�ͺ�@7<�&M�Q�6�
+�?���w	㝄-
���n`��Rb��[����]�v-��X�XXF����9Y f��x,�7Waʱ����Ae/h��P>;��8����C�%@U]���T���/���2*��1+#��A��zfp�1����(��= ��Av�:MKz�/x��F|��B�:ɲ:9<9�s�AX����B�z<�s#�sHb �`����Es�p!�+�[M��&���3�No� X�/��N��j9�V��Y��+aA�ġն���ϛ��{�M�^c1���_��M���)wLU�6ì�u�$:�w���y��"��1&�\	܋r�w���e̱���a�2�TŢ��r���Z��z�lZ6����I���2��"�������i��}W?����S}���I�iq��>�`�z}�����L��)�U;���4�Ҁ;�����������J�`]*����!�bk�T�>|�����/�PIw�Z'	}�#����C�HMރ01����blʃ����R�����&"���,�gU���%��c/\�J��11^jL���BW�Z�� <�޼�PO^+���+1�����@C�{��=�� a�d��
���jm�'����U޿{�&H0�G��J@��m���T�m�+���Պ���u�t���"۶���J2$��r�K�N���d�,������P0��kǚ�0֕FO̩|%��U�+/�WzoA�4l��UL��5)	�Mn*�LH���ʾ�C9� /�JK$���g ,w�K���v}�>T���+��yQ�	O��\��b�A 0��l�J׈G�����,)���A`5�F���F��$��]���ۢ�LE�E8�E[ˇ�����������ӸpF1�D��ݙ�G�b��JG�oa S����}�O
}d�(�>�h�WG��OT�Xi-_���pg���ϔn�ۮN�7ߤ
�bk���JH$������nz�B��{��C;t�y��{���8|�Ghrt:�3�3g�(ӕxM�T�>���vYwG��N��������4ї�xG�P��N�4C�c��)e[Z2s�R�T����zY�7���e�������[P����G�rɵt���-A`:�v�RC,Ep�-vj����P���k410r5�bq�P�ܽq�7iJ�q���,�H�m�[������e�o�:�_�"LMPAa"�����Ù��;�'� ���;�Kb���㳭���L��V�_�7�*��p�53<	G5�e�w]��& �@��������u���
����z3Yp�$�-����L��]�cHd/T۲����㐤�2�S
����+<�E*@C�N�⣓��
9��6;0��MRΗ^��lx����˝M�t������~]�`�S]��\ьC���I �� y��c��j�ꀙ:�@D�O�fN�|�s$���8�a��T�e5�*K�g���P��E)]�ċ{t�&W�<�d�o{Y��A�
�������v���RD��&�X�I��;�p��[�O�����Kj{6�����q���2=����A��c�� jB���Y�dfk��z�WO�XEAf~��^t�9���jY�1��v7�)�hOrl�U6�T�����O@�w౾�pm�c����wU���Amv�`h7��:v�^|�r�|%3��OF�/�(
N�q�}j`�EQ�I��������!4 c��;�SfviG7�NVϱPf&+q���L���}�Ꭓ���� �
�
�%>y3�.QvarE������[ܪ��W�6����Hk?�T��f������s�|�H����8}�"���°|u�V~&P��p<l��>��(:J��&�؁H;>�y÷?@���3����J[�!ω1�e"\���72s�MW�[,��QsK&�k���QV���<�&��1ہ�Q��Zr	��|�x�����t\7A�F0�+jbI9���5�|����P��03���ќO�?��P��~9i:l;�+���m�WbfYxJ���������R ��� ���܆r�܍5>Q��csAG����-�H15�˥*��x;E�2Q	q}�)2Y����ݰo�j�p8��ڊ���G�Z����k>WW��M��4DᦉR/�OP�g��<�k��L�'Cߏ�����7������Í�`����lP�����mR��O2��Z�ю:�'�%�/�J�~g���z�7�z�G&9_�M��<�iH����.()U� �R].�RY�v��4�<�ys�囊�S,p\�}�\�� ��-�O�����Hڊ~�zr���y��xc�������Y�<�d���c/KȨŕA#����H>1t� ��)�D5�R��(����4*	�Ag9�ƦMOy(G���M�h��7��yΖ���T��'�����`����f�lw�C�_7�r���"��m�}PLaH�c�����
��uJ�,�Sh�J�Z~ZM�r�G!�۟�{H�����Ɠ��L�ʵ`ar㆞�	ÄȤ�I�p�L`�`*��AW�N�
���R���T���8�q3#LXE?�qFΡ�{��sL����f@ȍԍ̨�{��NB��u�$4�' ���d�L �"��(C;�y@>��0 ,��/D��"c����=!1�����
}L��j�������H@���_��ᨂ�Q>�
r��7�t�X�N"dd��;�x�9��d����ţ��s�A��Pb����;�q?!���+b=|~���V��u�i�T�	V=^jI�A���E�gfIo�Aȴ�1F֮x
�;�E=�y�Xά ����1;G�8)�u2$��ҡ}�X����3����v#~C��G��^�m�\ tw �%��7�������*!2�߾>/ea�z�"?��P���]�%4ݐ��C�ç4�� ���M_���~�e ��u{B�!dnzA�����{��PY{>Vw�/��oI���?�����hFSn"u�'x/Ǉ�������	���אF��,Ǆ��o̽�a45�S��sB�����;�':���-��Ԟ�� �� �gJ���e�o��RV��dւR04rQ܄����年Y�[�Ũ$*�Z�ï�~�/�v������!������3��F�_:�_�I���Jc�X���F��&�o,��h�M��f�Dt(�_��Ԅ��T#�k�ih[hk�!z�O,�̱'3��Z��=M]��~�1�1HTZ��#�B�|���!�D��:T{�oV�v�f���W��~E .�=W���Ȫ�/��V�V���M��ܓ���[�<B���w���?�����x���C��e6P�cEa�N���]�v��j��T,����D���EӬz	���Ď�L�۫E�J=1Y|i ���7����IF��}!���f4���@��L9d����2<���Z���}�P���(j�lp�!�e�z+fStS(!`OV�}�c�q�:Ҽp����.!:|��n$C=l�|����1��ɥ��{��8g���1?���S�U���B lv�&����N5�������;H��|�`�s| ������(�B�&)�3=đd��q�)�'}�ѓZZa��(��&��S0���wn�(�ފhP��k����t1E�P��H$�5�Pi����6����.{u���7E��4r���{�P;~

�S8[	T������=����{�j�/t]���'��mB�h�Y&;�L���u������4o7D�s35I��_�- <���씥���� ��S1z�hT�[ڀ�AW��$�c�a �s�b�bvu B�g��P,ȸ=����������ق����*���y�1E?��4~f���aJ�h��cʬ�r���VN0���>+�7�@t�>*��Ia��>);��3�[BE���k�U0������, .���>�}W4:>���TI����ތ~h�PEv�����1@�ȶ��eF�_	��7�bT;��]�O�5���O�Q���9,��um�+ �g��(*�$�~�2�l��I�b���R�eocHx(E�C|�V:\�Q5������|$���-*	d+�ͤ#�%��[����u�e�?�2��ƪ%*�Ϫ�������F4��Ŏ���-��Q_w�?��w߂���)��{"�xՁ�^�����.k%����ɪ�aB�2~��h2�t-$�� m}���n�q+:���2�|��FAo ��K�Xq�	���R���a�T*>�wX�"CY(]J�Sx��y}�	�Cf��k��X@?X%��wؔ�za��� ���] 6n��b��T�<{5�~�\W�o0��[�4u�F�����g!V��H__F�T��C����ꋦh/�v@zGJ���4����Fş��ʑ%Rp%��Aܕ��P��F�3�P����������E+2(,�jڏ@p�;�V��gB]7�>�	`BH;Z��&D5C��IQ:|�(ln���h��#**�@��J�6Wc��sאC�-��GJ2���A�"7�CҢ�������O{#�6�t�.i�2����Z�/���O�4 ���C��0`��^�]Ŏn&~���Ʈ8��³�=WS��W7�R*���;���P��nMn����?wK�c��/H���4[��u3i�ڎ���(�bb�]�]>�6�y�Q�ރa+f����A��nn�f���jG������;c�࿶֋I�H?���z�Dej0��Y�Rq�=�b�\�{����>;�%kH��J9�'
�����@�D4�o��uEw�'2��|���;?Y��נd�;J���L{?i����v��
�ސ�+��Cb��y��U��5�M�x��� O�.�x��{�:��`�\����B����m����
>��ˬ@�N;>���+o�[L6�l�y���a�d�W[�cc��b�� � Z��Lv+�v>�c��o�iр*�w���o��s8�%�u��2jN �e:o|��F#�[�M��38�x��?��B��sS$�(���+��j_n7�5��#�Ør�����@6�"$(%�qU^Q��R���/����w�`��D)j6��^e5���z���� �|�t���g�|ې�䧕�Ƣ�D/�������1A�c&\�K��b��h�4���(_�i}��Ϣ�C	���ѥ# �[���Z��:�4�s7{%�1�l�ο,���Ft6���Vp�^��Ě���������0�0j��*$"��v�{� #*s��o>y���]�L�tB0x��8�F��҇���~�¨��]t��F;�;cj�&�h��jh�/"U8'�h7�����\yv������݇�=���s��0�S��R��"e�|��V��*.��'�b���T��ͤ����+i��^�BrN�Q�j4�����kc�%�F,b����#�S5x�aM�����5bF�0��`~m,�b1 o�SM�q�ii1��b6nN׍n�6��_�����Q#^������K-�k]a�9�H6:#A�5��PM)���(�%Xoy)����{����X	�f8�;\h�v:������߄[W�K�[��]����b9��@%�H�>"��}��y�)�
�*B�=G���uc�����*�J\�?g��/w�N��6�2�,��^LHV1ᎎK�C�6�(~Z�op���ȥ�n���G���yJ�nCH")�t_�1yd|n	�|�
GmP�#o��H�1|���ȝ� �wP��l7\�*We�J��L����.�z.���J�q��h��=�z�]���Z�������� f��>Lِ���V��<�������j�=��h�
7�~�W'�=���j�1;x�BqE�ϥ5�������v/�ďF��n��c����[�[ v*�5��mF]B�'s��r�������!A������ۥ��~�c��4����r��4=���ȋ�_w�u��2I���l����K(b�,e?�FuQ��\��,�3�Kh{�#��������"���g8�'�pR��U`�p�E���y��S�:�����D���/`���v������W�2��b�<�`�eW�v%��sկ���[�%Wg��_o�o���p��w�t(��6�%+,q�_��#8��K�@���}ʌ}���3���l��jr|r�ҔT<c�U�X��6'��e�<oi	��8D;
��5�J��P��'x�{�V��l���8Y�j�ݟkk�I��1ic�'�ߊ�N���Bl"�>�+�ބ+Q�~2��:!�J�\v��L0M�.$[Czs���4�v����:`�6̜�i���z�r�j�bB���3�>���ȥ8Qi$��&�|�3�r��Řk����i��G#*64FG�cXV����e*! p���J������q���%ᠪ�?�W��>L�7f�Q�3l¨�}�m����(��;��۞�[_��ϑ�u�&�)�FT�0�)4�W�a���"�)+_��|����4��
k�q��L�^�-�ޘU�Z��tm���f�]ܠ@y+r����j;��k�}�.Z��	�j[�gٱ�V����m4�X�!Y����f���a�>��D|�s��CWڮ)�X�������*{�mxH."^c*uj#>��^�ۡdM]�t�h��i2����l�$b3$$b���d�J��X-:�΢�� !o7���4���R<��*T����	Sky})�ƨ����E̬rI�=YP����ݶ!�iw�˵`�E�-�z~�#��\�4������|�����=����b��=�1����E��ues|wJ�Jm&����c��̔0��� ��	|�ľ��)B�+���h^ĩ�3S`��oF���u��t�6Wl��/������4���)��o?T�ta|3��
��[�7&��Ə�O��ȂG����],7�����O��TR�7�Tg<CL{�w�0�sk�ӏ��U~��F²5[���l-�U���^��%��;-�j�?���7ޠ��|s��ʒ;�BDA��������^/�?7Fݞb���Ų���e��L�y�:�q�|�|p�x>����1	��jo���M}��_M�-wF�Yb�I�kP��,/�!���V]��q�����#�E�����f'�y�;�.OA��6,H�=��;AGI���X�z<���W��-��=�W�""�L�i,<Nw7=ASamC�(0�Pjr҇~�����ӥw�O�	����&'7<�;0N�X����d�ȕ|�n|����2M�p��e1A��uwB�*3��OW���EswvW]��"�m�����Ģ�Wʘ��d\�lQ��k����X�B~>�y�K�P^��^�Ez�!��T��19��Cv<��(#�%Լnm��9������j���?�4JЁ���V�.��5A��uF}x{d�ӾAfJB�R�-9��>�Ä��~w�o����Nb��%�?�,��Y����<c[M���[�!�NY�a{���G�l�?j�L/�xM��d��6��[�M����_��'A�l���w���u-Ҷ[צS����м���st�e:���	䍺-5i5�F�6�쟗���]�9�u���,�����C/�,�����"��k�u�Y�"Ǎa*8�T	
�h>M�O�1f~Y��4�a���fWD�)� �2�3�XG�>f^�ۯkp���Ţa��r�N0庝�d�r��K[ɢ�y�����,i�s�M��#w�耘���J�|�pB�_���~%�/���h5�������-�O
�U�����ʳ��r�a��o�>��[��@u�n�� �X�.'�*bӼ�nlt��x�PI��Iޓ}�݃\�Z�j�7>w�M5�7I��/�ꉪ�_��R%��Ϲ=�QK�V�T�����;f�?����+�eg�Ŗƾ���|Ì��eG����]��b������J�&$��˝����֥@݇���6�?Sn^�ϖխn����^e6uz��QB�\���MJ���yϰ��r�]�۳��
��+Go/C���&q��Ǉ�҅�����<�"7��P�ϫ� �)��{L̲V$h�Hk�O޷���S��V���am�V�5�g���n�i�*�}�0&���Q��O�J#s�����)i
����\�]����ݳ&i�ӄ"P���ũw{�`X�p~�6j��`�HT��O:W�0q�}r�O��"����9���8ゼ,�_T��"}�p�
��Vl��#w���_
[,Mc��wJ�P94
� �_����)�p3�E}��t~B���9��u1�Wי�0�J̑�ZH���<��_��E�x۹�G	}��hq�h
{<c/H�͌Y]�D-vGYor��H[���mO=շ�"}�'�5��>N>b{�v��^�zMd(t�^�|=��&����:`�����	�R�.V����������;���y4�Z�q]�)c�^�:�k�^w�Y�~6l�~���~ ����I��ۂ���꓾�e�֕sPZ���Yr����v���Mx��nSCG/tN�ّ�Bm�Y���o�\Tj*
ߑ�P��|�������}>fGj��R��MMؙ��&�u8{��w'a�����_Kfb�DB�'�]��ZBto�%�j�����OƦ� U�c.[w����d��I���^D^�W�����nyy�#�*���&����+�ȏ�c*7�З+���B�f�ob��0y/�k��� �fأy�E�K��Ud~��@���"F��%-�K&��\N=24�T�P!��?ɒ��B��$]M�w�S�4�,l�� �Eq/�z��~%s{��\��-�y�-�.�{/�z�oY�c�,c7m϶�s�J��Qf�U�toa�Զ*|��� %�v$l�Y��Vހ��Pe�Z��}�1T��]�8�!<6m("��ͤٽ�}�9�i sY �Z���܍�-;4�^�?�͛��Eq6܍w�7�,U%�{&-.>y/[�oo���u��M�xYJ)M�Q[�AL@z���aI�NTR���J�D�A*��+��7޷}�&V��g��3v��cL{���cNc��5Z�vS屭������? -�(6��%�0Õ�*��`8��%bVR�u=����R�qU��~��v!� ����U�&s�9��	��}�)f�2sW�0�U43U�C�ޟ.�=0B^. <�ND��c_މEb�"a:򨯂�\&��qr��Pv�FZ�쬖,�'��/�� �3�yv�5kL2r�[��5�����k���x>�}?���r>�X�N�Lg�^�>J�X���5�";u��W������l�:d�;����<{<�^���c�s�'DA-1f���~��3��C�峍����qo���0G�C�z�'���;"������Q��n�A]���߷����ú��������	���JI�mQ]����޶�C��R�o�] �G�ʞt~�$��$���x��?NC?��@����
ǺDN��R�7E��EkǄ(C��ͩa�,�1�2��|e�u��I�����7��U�]٭>%r�/�x�djO�-�+�O�mg��x�<�*U��1�=_늦:�^
����KL��LH]�L�'l8���V�S.�(f���ge�N�A
�!�_����S=^
��*|0؎P��	���uU�Ƈ�锉+H=(,�0����A�şԟ�۟S=N2?�{͞�\5^_�97��K\IH����2�,Hψ꧲b3�e��ݤ��<�nʛlҟ����K؎�b��*Y�3Ǭf���<<Y(�,�8<ۖ�\�-W[/�\�X��=럯��4�>?>t.� �`�4�	^�Kon�mX�]\$��Y$�?�n˩�k>��~$��~�p$��>���gWr�*u�2�6�d��,:���9�C���\B�й33��5�v~8J���}�����ؖa�>�.o�o��X��<|#M,�h�B�i�d���������%m^���ʦ/�!�A�'��dL��J�t����I�!vV����`&ܺ��)�s%�}�b>[�/��1�>d/)(��R\*�d~��?���)?un�<�-X�۷�<�(V�U�ˢ_�&z{�ʻ�W@�<��H֒��<t?�h�I�G��ar��L����A����Jd]���O���+�MQG��Ke���ZAQ�J��^�W����֏�������OM�G%��֛u��������.�S�����&
#V�W-��V�e����;���>,�Ώ�;�{�o�����Z+~dO\�J;/w�����8!�6W��.�F.��U���k[��i�`6���Y��
�ģ�>�p�^ta�^  Kr�bG�0�1]��i;|���o�����y��voTm�_���=^=�XvS��%fJ���co�C|\4�{�e��/<'8m�{���j�^i�~;�8���v�xT���k̃��3[��ǭ��Nm���w�������S\�P�x�ʾ}s^`��|^����Wن���>bd�����THz|�v�P�:�&�U�f�*��E#�a��δ��G��᝱�(��4��
���{g��M��u-����M���ֆt�}y��n[����m�$�9G"��K�ˎo[��7sɛ�:���{X-��.;�/$�l���oq�W�x���`�(���V�]O��|�ޡ��Z������~p�t��t�#}e'�\u?>���QVGQ1�|dR��yxD�px}Wwt��{����	k\�W$�N���wM.pބG��~���m�+ �מ�x�9���؍;<�6Oc*����}�
O��UfR��Q2��jR���Z��Pox�=���1�*��Y���p]�y�����/��i<��\ŗ��Wx�Z�X��pg0a%�~�5�9���T~KN�y{}���$���8|�Ik� �>�'��Ey��Y��AL��N%$�Η��Þ%�a����Hd�m2lCt�L㾪��~�I�Z�?j2��d�ݺ��1�^t�ӽ�3>�&�ڙұ!��j�b۟I���:Vx�������u;��xl ]�[�����oW�8�gԥ�w �7��L?^vg4��,O?�f��"_ٷyw�/��x�>3Kj�0�m��la��eA���a�8�E��:��ʶ��Ƚ�G��q�삥~�ӯF������A<��L!R���Go5M��g�]�)������q9Z�|C�I��E�O�G2�+��o˛�ĳqj�a�����D��m:��F��&s>@*�~Ͱָ�~Y?�<&>=ܞ�l��eɮ�O(�ٷ�P��/�d��E�O(��0�qj�-�T��޳�EQ�wִ������$z��|���c���
_{բ2�$q{=�de	�*�B3R��k.	毓�~'N��r��WvH=;�<O?_O��r�%�|��U ����5�t���E��es�^��5�C���G��L��A�ͮ����YXq;�?>hY�{�`	�!�t�47�/t����\��V����о����lD����y�!N��+|)��Sг���ls�������|��������f�{���r�n�#U�樹�)�#1O*���/Ԥ�LȭA9G�k���v�?�4�ɖ�n�#_d�ޥ7��K�<c���
�)������ngG�h7���,`���d�,��7��oeD��cE�@FU0�wVm$��5����h��о�.B{���nh��V��䇹���.������@Hj��� ���"��M�N�cELC��Y&E�A����`�Pm�.��G<�k��	Q�ͳ맅[�u�(M��<ߜ;����i���߬�n����2�#x.����ɝ{������#�=�jV�u�,�.M/�<ȝ2�����]�;Jy����{�ط�:2]�Y�{�b�����ݧ5����.�n�~Z�|�/]��!}��U{��k����e;��S�#��J:H��L>C=�/[� ��7
/E�s�V! =^jY썡^,Ѭ^H�sXHf7X@g�݂r���������
5�V4Oa�F8����u��ډ��=`c��U�T�,_�A���^��D~�I����އQ%w�|ӷ�J�Yq�+{�d�U���mX˻�4��,r�4\ ������8}�+�)��6�C\�^�e��w	-k�g�����/4���*��|*������^X�B{��>i��p�a<h�ꡰ?�;������1��yٻ7�����vۦ�rJ�>�m�([�fō/!G�>_4����x<c���6,�n�v��HZˋ�����{����qS���C������ȡ������ �շ������Eo����Y��?Bֲ�j}�dmT~&��������r�P0|�ګx�0"xN"���6q^�p��s4gQ>����a�Snz�1�+]�N�'B�,81�LA�ai���c��_����kOL���f��!�b]�U�y��˚S�g<dtu�
�ŵ�11�D�-�6����	8���U�J��c��ί��JH��>$�@�S_Q\;k8��Vp�ni���h,�+Ğ���WF�q��0WEVV��Fg�3�͢ÈP���W;"s�K�޷]�Y�Ds�f��=߬GexqM���(U"5�~���梗�/�ƶ�h���!�˸��Y xގ�/�趺*i��x;�ײګ�yb:B�ު�|��7���W�{�V\��>A�N�n�HPjy�_(9���{��n>�~�����赲W���eo�eyh-�O{�n���(�g��J�(��w��VGg~��7&q���0�X_�ҮP����v��E~�`Xq�_�U��Ҭd:h�O_�)H���]
\��Z��S�ґ�Ud=����V"}���K�T�s� 0�W�yU]X�'X9��Mg"ҙG�1;T6�ߦ,0������o�:�"�Ww�? ���}���`P�6��Ԅ�,���s����IQ��2I526��1.��[ӊ�y�ϫ*���e�a���>�vi65��������f�S�UebH�9Q���kq$�#D���a��s��
�9�{Up��qW�"�Hm����3�������B��y����{��`ï� ?�(P�26b�S�̟5�"�i�J&���%,p�cj����E�l�1{C��OI[�۶\8��%�9�����VeP�P��/�_Ϻ/ĺV���h4±��T+r���9a���Ԣd����a������D���za����|a	U��^�`���VLU$��|A�D�r����'2�AT��E�\��l����x�,?&r��eٳ�}-�^�봋`������~��bc�ĺa�Q��љ^iݘ�<
��W��HE�)]�k\�W��n�����U$r{����WI�l =&*5E��8zi�GH�R�e�i6����������k�2au�]t�v�!}ft�
�*"�\����j;J-b/���m�(�E^�_8�ځ��B��Ù,S��?���E���Շ�$�鯞n+���n��l7�	e{`�}�eҩ>�&�U���6D���y��qjbm��qI��+��|p��;y�-,��^$�2��Q����|�QSSο�˚�WǕD��)�ɸvE���Z�����3^+�J8�a�U���9k*ģ���"��_�΍�w-s%���kd+	�Z�rM��
9�K ���E�ǔ'��~��:z���E�R�Gr��;!u=�yZb�g�I8`u��s7fQ?7��7tR�UI'�Imt$��V�?@�5@i������?���ȏ=1n@�FS����_?�Q�W�|���Axڛ��-���C�#ܲZ+���X4�h��u��V��PH7/ƕ\�E*�g��$�z���_��O�z� �e���I8"PIڠ8^�m�f�m��qг��Gz�e������� �6��L�GO���'�)���W���
 �+��q!H����C�YE�6c��V=`��$�1c�l�(�:	��K��'0�������R��/5�l�f -�a��ᛚ.�'����%rFe�2�/����?m�E�c�`8�	�ַ�!˖mj
�� z�©o�he���7����wV/�UC���T2�M�ϭ�}�qF�.����\��ah}��+%U:�x��0��(t����y9i!�֕�DW��b�`�yު\��+��?	�� 1Q;)l<�f�'����v�"<���V�G(��ɲc�hy$Ԯ�*�I��<���h���$�T��H�*��-d{F+��q�%�0Q�� ݌�ع�`#��"v*�R�u"`�W���<�ڋ��B��<P��vϸ�f'�JD���,':p�bu�>=�����c������e,�"��Dp��F��S���\(��AYL/8��*�:K�u�_g/\�,_��@�$��m�_g�_�=����R��~��N�9���3��pZV����P�/0�׊F����F:ylQ
w~	Eum\�H����'�3qW��/���@=W���1��og1ǳ�za�UՁZ��qL)�+�d�9�ǆ�@����4?�}T� ho"Bd|��j�B��N:�n,��-�E[��7otl���;)	��uT�qOS�tp�qT��,�}���9�ְ��-�K@OU��}x���L�bki��@��sԸM6��~|��ܷ�g�+wIȞ㤰��tց%`��@]����L�u�@KJ��t��͑�pq�KB��x Q�����u MG������d�7D}��A�3�`С,�����[�	��
/C������"�R�ҭ]_��G2�/���kvj���is��9 �  &��gb� ��]X�IdC�U����t���17���[�D����;y%0��A����k���3�)]�Ō��U�u5�y�1֖�1�(����Վ �W;����ص���Ҁ��Z�i|���v�H�.���O9����Md���\��`� Q�U�
�g+��X����[L�3�b,d���W�ab������U�;�6;�_:�UQ &+�f�Ct�X��T�Sk��Yx����EV[?�J��o+v���php����L�'m�k��W�����S~�@�^QEf�b��4JTe�փz�C����y>��W���c&��Q�v���Fmxy��+~�eYj��� �>��b0G6�����#$���F��,ZH�
�"6ї�<��S��эk�LFI�C"��b�w3~���,��W�۲���ׅt�p,.4:,ޜ�W��V�����u����V*D.����HH�U�:uO�䬔w�gViL~P�1+��q��|�Z�_jF@Ly�'UV�\��������e��K�ض3���;�29%t�o��э�x���ٱ���ab�v���8=��27߱gh�_�I!.�`9K&+<���٦�Gc��O��h�kܚ�RO�Qz�A_[6o3_�y�|DĻ�H7C�s�p��r/��M�&��j��$l�T H�	��R��#s���Xm��u����#�lTI�f�����C� ��-Z�J�Uʻ�aXw��]�a�m( 3*��V��m����'`)��G��U�倸~BW�BkX[�@9��@9)
g0�ӟ�u�ǰ��W�w2�q��	&Dm���An�;x(x ��i�d�/�*�Bd�U �nt�Qڐ����U��7	�:������Ŏ$ᱞ����RJm6�i[���j�7Q�9�[s�r�Y�p�jg��l�d����?��������r-��<��9ɩm9mеUT!]Uؑ����(��٭�Y	Y6�ym�5=XK�^��xlHe�:ʇ�B6�I���#�����vD옕4��M��5�65���UZ-[���]��	�UjSU��j�ZEͶF�7��?�s��y>�>�8�9'T|��j��6*4gWi�yl��T���L�{Mx6֦��h�7�AbƓ)�	fd7��E�u��
_qS�BT�|����S�#㉺!��Oo-�)(�TCwJI��ƹپ�g��]�hv/�zޒ����h��vZ��:G����lR2@�/F/5];��?h�yۮ�\\��;��߹�ut��F-4~!���z%,(�CW��t\���A��H�|�z;K�3����Z���0��:b|�����������̱w�]���0@�J�L"��R%������2F�Q���xN��	�;�$C)>����"����tM�F>�DNcB�'�NsC�>�R�ngrf^=$[(�v��z��饍v��������7�}sm@�E��f��rN��$G�$�=���}�[MYīprlB��W�{x�Y�z_���D�����s�Gl����_�ЛJk��DՋ��D��|��`�r��y�j���{^����R�!��]�Lx�n��52C��Q%��_�Iv�мz��[3S�K����&�\1�S��(�r4�W`���9T�T�c���[}���S��^c�,�zn !jq�!���F9��Ձ�Ȫ!Z�, ��p�`����L5�2?,�e�����M> C��U�[/;3���xe"`U����E�d6ebA��^P��C޾���o/���J�Lȧw�a�@Rn�b�XVݫ�*��;T��S�м[-�Ow�UO��T��h�l5ި*��JiA8y�k�S��Y�S(��Ze�N����K�ݑ_W����.9d��2/�=-��?Y����x,����弗���Y�>bF��@��L���#�kK�$�4�Kb��+_;�A,.�苅��NrT$N=$6��vϾc���&\��j-��wO���,���L��G��ӽ��ÕrR��KH�����G6������C�|��@X�9��!q�XyQ���c��;��f�|유2OdN��gOW�WX���t��*ڢ�ı��xx�3
N�����'�p	L�w?ɓ��1j ��G�Rk��RG�νO��U���|Sg����N�Euִj%��8��_�0u�,XW[eYbT��%J��ۋ��{���D��a:]Z�����l.Y�1�%z˃�#ۚ��,���Y)�<&�G?�;2��� ��3^����H�����\�#�vsd/���x)�=k�u� ���I�=�q�#�J^.�������r�h�N��Y��K�&?��F��\,�)S�#�@^ ?����q�^~�J����l:I2��Z���T�e�˫��7�_?��<�^0����7
���N��P��4��g�7]�ǥ�֫
���];h�K�Y|�q�t�{rE����&��e��,��3����wd�O�X��Ч�e�Ip�OPbm�,r� b@18�^ᮩ��[;1��߳����v�^��A��w�(�<|�٣�e�J��O9�H(jg>~D����cuq�[���$��|�magp���'�"�<���(�p}���{\�@����1��fvB�t\o��,%e�!&��YeC�湾� ��A�p������y}�7�1���	�h��h�<w%*-SX��i�h��x���)��#jg,G�;�"��kdQ�6�h +���-U-˜+V��e�j���}ٿ*��p�n�y���%R�؅<�y� ��^��"�5���b*X_~z:���SU���?ƭ������Wil��8������I��\���5җ1��xk���{�ٗP�<`b��E_�O�ǧZ|6�&ƚv jZ�ğ;"�e�N�;�VOL�˷��?�]"Hj�h>�]V����<�i�qo&,&�}�]Q6�pU��`�@�T�\�p���b*�U�����E[�:�L�排�����[k@����|1�4xq��3���_V��2�u\�A�b�Ƃ*�Gm����5��DɇQ���G�?����*�?3����!7X�����t�������u�خ#Q��K��	u��ѣ��:СO�̋w=�Cofs`MI؄�9p?�P�ޏ��I����#���{�gJsl���'g~�����<�B*Oۄ��������OB�1z{�]8�����]T�Zo\�C	,���
�8az+)B���H�ŋ�~�ZI��)�}2=ބ.�s�~ �N�ì[�"��oUx0]4ʧ����2�2/0|�#=��J*�L��l+������e�$muV�޲�n�c22#�[���Q���j %�@M�Mt/��z��.�OAНF<�T<Ͳ���W{�2y�}$A�����<��W��m7g�G����b`n~=u�kR��8��U�g�*���Q5���[�3"B���R H����ڑ���@��H�Z{S���֧��~����9�B��czw�Ќ�ԇz��m�:I���I;����w1u�t�u��˫ƌb�jŒ����a��4��T �*P��^�#����ҥt�jL$����*B�����5-�^��xZu(�e�х�6C�����}'��:bV����K�v�)6ZV��3��|Hq#l��3\wȑ=�t"�j��л���zk���;�||Yxj.T��+��/����~>~*)?������f�
�ǟi{�G�慷�2�V�Y�<�,�34��A�)��C
Ǔ :��3�A:3+E�b�a&��*k����v����&�h$������rr�n>>I��[�7K��՝���)M����@��"J����|������6e|i��>a����Ziu��=����K��$12܀정V���V�}lW�\�0�\k�'t�I��!�X���ƶ��o�9B,7�`�� �H���rhŻ����2������gB��V#����Y�����}��i1$�ֻ���|� P0q,�z�rV�5��A&2���J�r'��֪KU��t{��H�c*��<h��`~^��go%��j(I�>��Oۉ1e"Qb-�W�^o~]lË��Ľ�7��h���!wZ>��\?�,c��X�B��uI����5`�^�i�L�ʫ�ݱ�������~T���~��.���g�$	��Sw�p��+!�B��&(A����d�F�Sᢱl.�DJ��r�M_4���Wͩ䎻Z(�̼k��'�
i��4���J+J~�1oQ��r}r9��/���t3�PV�Đ�p�nz���[�a�V���RF�'ai?Y8 a�W��RK� @g�%-6�AT��������M<�~QY����R��m���SVd~����|POX�?b�Q���R�0�MB���C��q6���/���P6����FqB�}Y;�Ⱥ|���W�p�L%����l8�ԣ�r¡6́T���6����d�~���C�Z��P��$O*n#����	��O;�H�Qf�W�=��=a݋B�=$!�Շz�]�O�SAjr&�M���'�"`��_�E�O��.$"�2٨)�}]��BQ�-�u�����ܗ�:������S?.�(ZG�G��P-�m���
h+�Η��SLN�{�	�s8G�]���pC��&��p�S����hc�d@U\8�u�Q�]��7F�'�V5�����������/Β�O���������p�b�@��`-V|���z�P�����k*�H��.�5;�jq"�7�i4�z�d��t�K��w�.��y�fz�gq�yƸ��b��=�:D@���s��n�ϐ��<���
=�\�.�줻�La�;��T�h�\	Y�`Am6J:�䗂���!M�k�$g�� D�SU@j�\��"�7S��r�r9x0�׀29R���b�h�N��%ޖ�l�O�/�%�E�'���?Dn���L�g� ����NE����c�@	QO��Q��ϒ�za_N�@aE~&z�.Dg���i&�ou�����X���D=�6�rWG1��=X��vGԩ]���A3�Z�����b:��I����L8x����9��=����.��0�����������T�,�1��za=�#�9��}nv�C�̻ܠ�ٸ���S���2�d�����Q*�B@�CSM��|��$���"z�n;��W�@a�8�z��Q����>��� �R�����cŪ���9�W���b��bC��I�wɟ_Ɂ�U>���~�}�f0S��3�����?`���G5�<�qȅ��uX|8�r�.1�P!�]��[����f/�,?#j2
��/�G\�����1LĒv�~.�)���ޤ+�<�> �d�X�I��"�]o��L�Jc㖗%]�s/;�T�y �WG�p{�,��it{�s9��P|����[���i@�Q>�B	��\&��Kb��k+��'������d.�����8��;��e�2a�h>-J(���,����'�4B��A���C��xE�Q`�h ��l�k��7Qb�Od�瞷���~���ħ>���[��>U膥rA�0��cI!سV�
I�l[Bw�^"��S3s�".�9p��n(<�3n�g9���<.��MC��}�X�j]=Bjʘ�r$ĤA��B*���m�AO��`�JV�}ˀ���gA�� ����1���l��Q�:z�{�E��4�� �INŌ��'�V{�]��4U(�2��yِ=���u�-Q:FM�3��[�ݨ1׊ܿbm�(��&:&<J�צE^�B�0g)���6��V^��@kY4��E1��d�?��o�4Z�2�}�m�Ld�z�.���Y���#�&��r�W,�׋5�ц����L%E���n�Y�}�t��VeB��|J2�R���²��m�r��|6��߄�iX��j�LS�x�eAO��1Ҿ�0�I�QtoA&<��� %"$�� 2}	��PT跥�Z.��哯S��=�t���ט�����#|��+o�@�j������Kx��+�V5/�t���^�-ar�3ʛB6�-}
��a�$IK�ې[�bY��އbQϴT(�_]+�M�&�����H�X�{ [��LΎ`������P\	_ي�J�Dd��&
��뗋�mc�Z'
�RnD����a��"~tUS"}s7��bw[R���|������'��e�*���RV�bP��p)�W6�삷1-۸�跦�h	��:���רÔ��ֱAؑа@���GtM{����]��Pm����,4�4��x���JB�a+�������:��L(�SH=��_��%���S�x^���st�O�����!��,
���aM�ϛ%�VR�^	 �`B��1�$�J�p`�H�Ϥ�_���	Q��������c��;S'� �M����q�U���K�����ﵹs����g!�-�>Ŋi��Я��B���X�MY��1RQ�oj�-s�Z2-���"���6��t�u���:=z�-4�C@�t�]�YK��0�
���fP�ē�Tv��*�����uؒ�̐Ŕ�}C{`��:T�ɵO����u3�!��Ux$��)7���9`u�VyIg�s��h�L(ܜ�ö�R0 ,���������m�ͩ��ǐ�U�	-:��[?��`��S��y�>'�|f����e�t-�&�8]slp����X�T��L��DWL)���I2���u��H}�"B_��0�Oż���0 ��jw6a��!�c%�mh�<"��>�Rp�3�C�V�4�����ǅ1&��_��섐]��U����Zo��N��Y?4�p¤�F+59�U@���7Ӥ�*
�;�""���P*�����? �z�h$�� 
�Q2$�[��o�o�%�Q��E(���QM��h���T%���K���.��;�lU�o����7M��O�À<#������:��7���w��x��T��'�Y�"szb��/7Y�T� Л�5'��|�� �i^w�r�DSL啍I�qz4�����i��CFMl)��|&�րZ�z� ���}i{��*��?:\\�����Sx�:/k���g9�t��P٢���lO=:�S�<a��9|�׽��?���''���&��:[��
;����9Yv�/ #�J�/��ɁMF̩�|0��hS2P �,�I�����#�ds5�-��RA�z�&�y�Uʕ�쫙9�%AA?ԨJ?{^:"�1���P:�BW�	V?�(/�v~#��G���"v)[{BIN�3�y�����Y�=�^/�{���^eS|mt���s�(�#�r(��O�^�Pj7�D�S0a���po��1[��\�mO����Ti�C��́��'t��UJ�(�cO|g��p�R4"�U�����HQQ�#�xv"�Vb\B�{Y3U��a�s���E
V�l���ukC�V�8]>V�}ߖ�Ƿ���x��3n��L���߀��rh��b;Ъ�O��a��cZ8��c��RQ�t�����m�W�Qצ;�B�B��_�cSN��͜
-�Ep�ީ���9X�tw;ȅ��#"������i��.��I�m ����Q���Vv����)c�osd���b�*[#BV�f�l��;{�&����]5����+O�!��~��6��6Q���|UU$ա[M��P��DɩU�P{�P����Q����C�.Z6܂��@�����m����Jsj*����q�� H�0�����의�˭t��3�-��,iX������Y����#�
Ɠ3�=��{��/L�g�г�J����״�a-��x�'mW�u^[xT�ϗ�c�c*��ZD�PXe����KW��z��{�1��Q�������hSY0OS'ਲG-&�ױsD�Ȥ���Z�3�߳���n�O�h�ag�� �=�Ce0}��+�s( OЄ�2}�|��(P��"
�-G�Zӕ���/X�-�>�p��}���dB��k�I�Im�J���m�ʈ����J����6�an�P��jg$�R����Z����3�~��"��ׅgU���Ӓ���
*l�2�*x�Q���j�������k�7B�����"1���w������K��3�����Մ8��!+|��´�0��z�i*`���rrd�́�/&�HϴF�EH7*O
�/P^�g�*��ow�v�F�,��|��i�uH4�Q0�|�Q�h���5+v����{e�E�뷼/8�T��s����STUY��C1�K.����!��r��Ch2+eRA��곏{�	�"��|,!kE]��#��ɹ���[��y3��&���}�y�j��|dj^���� ��>��o.�[,�@e��[>�_��;���⧎_�J?�:�����,$�};D��!�i���D)����p6�tq����S=���o��u�z���}���߰d��맬&��r�d�:&��1���c.勉�]Q��P����%����f��k��Ő�
�:��а���n���ķ?c�vL?��X����F�����vQr�a:w(G}@��~�Z;�
Oe�WH%H[��ٛ���,0z]����e4���z�d��="*�����v� 7ب!��Z�-+]kC��q{}.��o�#̘R��yF�`�TŰ��0^�0�t��'��/6��?W��`3����׏�0�#���Z�^$�Z�3���qG$�aqv��GprE�6j;��7״K����U�$;�.�Ym�Aiyl!�H��
�K_�nH�ú����ʿ%J+\]�&�h��@C�ű�$�JY�eY�΄�V��ܜ�vO�����c���<��q�H�:�t���6Vo����_��eW�,�!��?��D�9��Ā5jd��,����EF��w����۸H��u�s�֚���7�F��b��{�\��u�T������٫��hp��W�OKv���6��0�D�ͳ�D��&9�dq8�Q���qG�D�r@�B߈�8�i\vC�)
�0O�%�@�C�F|q�G?6�3���Eb�)�VH�/�+S_'K[F�9���J����EJ7O"�o����#t�ٴ�l��ޯ�ku��*�CH'��M�T$��V7";��e��n�^Z�g����o�f��vP����� _�����]v��ME�	Z7 ���W���ĭ,d�P��I
%р�[��~���hAO��^p�5�,�8����m�r��J����!�#I�Zr\�=���,<�*�3!(�5�n�N9*g�<w+S�n�V`8��r�빆�aўS�m�A>�h�A:��唦�#�>���2V5�VZ�]:��[��G�0�U�c�BIq#&[V����h}r�kkԎӆQ���Q,G��:	�ZE�ձw��Y���1p���4�g�N��pF���|�YhY�Y=X����Xx������!���{��C��m�8e���HTY�d�ڲ�w�����+�Ų�� # n�޷��̦yɌ�"F�cZ9M�MUq�8��x#�<}�����p�ua��z�)Z��(+��OJ���v��vie���Q3�
��������5�B�V7�N�V4&I$���4!_���o���Aŧ���9�����[N���"(R��S�f�∾�?��<��jQf`b���/!����:�֗� <��u��rTCA^�Mb�||�mת�$�S���m*�W�wNP���&�����WAV��������k#�N��@����uY��E�h���Z���{�l����ɝ��S�?f2��y�������ã��l� ��+��Xvd�_J,,�[�*xj���O��)?!�*�-Ja�G�Mu��=r��V9�L�b*%B��H���7��e8��_�d9�i���O�����&Do��|<�iq��f3f!����;MY��������	�����|Qb`�d�G_���4Ʈ��wNH1v��m���$��y��m#)W�x��]�Q�h$I�C�� ��ˊ��C�&��l�Ni�V�H5[A[�,7���<�({���K�?�f�BI{�}tv m�A0���42����f+�/�~M�,� Ic��`Qe"�GOu"�*G�	N*Rw�IP��|�2d���8 �{�%�+�I��_疢�̀v���ֱ����	�@zEŌl�]몢eE^&GX%B�Z|��l���l�"�����)a�xcC����J(k���:���v���{b$��u�wB՘�U6&u�e{�/��&�_7 i̓�cp� �.�7���9����|�X�(�`��m�t���Cl���A�߭{�F�#�:��X�y4��2�ww�n�d����)���}������1̑��^;}>}�EXT#�E�,Z�FTd[׍-����W�;@�CT�!���Ȫ�������'<a,�3�[�q�6�(d��).�q��Xջ��l��~/���e!3}�EJ<I��}@"5�&��I0-�Q��5I�+�;�N�(��{�Zy<�3�WT&;�v0��ԟ��e�p:f
g�`�U�����h���Z ]���Ki=o3p�IF}�>N0�rӠRWr�Ӑ�\*�)���܉}>�zgM�6|O����̿/rN�S�f<ץ��W��U;�ټilLǎq�v�A����\��E�X��eDr��ǅ��X�jP�$U�+t� ڝp10\ۘ��E�8��jx]v}�h�E��%�95�Ib9��_]��ilznЎP�V�(�0b�T-����=�g��z_������b�o��S��V��C-48s �����1h�N����%s`��O�᫮s��<m9X��r���j�0���� �.�Z.;O1rc�G�y��a��!7k��b�h�Y�_�+��6��pnx�Hgo�3!zWX���9b�/BP����R�-�
���M� ���mK�\�~k�W���D��k}��pr������u{u�R6�h�e���y2�J�.w�\k7*��O��O-]�NŪ��A����j'��!߁N��]��05�T���� +��_=1V������pE�|���2��_�"-�T�k�ҡCd&��	p�v�&-�??8��iHs)0�[���@��r�u�^����P���5BtHߞ�I��kGa����9�&�u���ۑ�)�}���vp�p>�!��C C@��j-�WZv愠2�-+C��Xxi]�T@�u"Jԁw-��L	�шqG��L����^��ԥT��ūn�7j�<=�ZizF���[�[.��5��j�|f!~��Je�O�ɟ�'=�1�Rs���d
��0�������SVv%%>��l��8��Rz5�?�Bb����T�#6�I�R��^�&�!pC�C�,����w(~,��L�{����g��c�������W'���Y�9I���o�!�����������gm���Ղ��O ߬��Ruj�w���;�Ӕ��L[gd�J;Q��񴢛����|>��';:���Ӆ��~!�<��>��]A+�޾�N/2�I=�Hor`�>�����/�Ŏ�2(�d"A]�F�jR��{��NE�H@d�w��B��8��m+lt��:���-$R��$�:��YI�p����5��zc͗�eÔ}F�t�_[���W��t��_Ϩƭ����{R���3Q~�=hO�_��K.�!�����v�Q��q���ɩ�e�8�j[����^�������B�?� �� .��/ڰ�a����yS��&s#ͣ[�U��fv�M�_"�<G�W&��#�Znq��˯�7C!)xD��<d�uf���Zy��R�����{f�n�}Q�s�}�@nfύ��'d՗W}��\�F*�r���C�}�TF��bEٶ���=6�{8�x5sg�.p�=�P��@����쵃���)�FC����ۇ\��u��S��[��/�{{������%y�(�B>:N�>E� �>~�i���a�&�<���۵)�n��,Si)2s2����l0��S�B���X�Ķ���Ļ0��7���|����X/*r�q����&1������,nu�<d.^�ق)���m=k�&]�lH��r�*̭a���(�i4�6~e�7mci�Ik�C�4�V����8zH$�G��O9��H�hO���3[J����^��@�X۝�Y�!� �ߡ��fƻ�>�A1`΃��L�j����%T��=˱����K���T��1s���?���s_���Z?��Z�����^��=D�s�@�$�R�co%D�������&�}�>6�N�7TfY<�Q�Y��;����9S������.iO4������e,�}�Չv�ǵS]����(�h��K:;���z�c{�I�_p'��,&��8c��C�����S����
�h9kg/I�	,ce;ؗ�vT�A��;L���r+ImK��?�"�,�1J�漞y<�q�cx/%���i���S���y����^�]�L�S��<�I�����k������к���۴��h�(K�-K#�$�+�Ǣ�^�N��L@��]녙tc�����b%�-"�Y�73�Q�X*Qg%�1��y,w�<ˁ܌���������J�rd�k��͈�[�2�5H�q|�Di?�l@�T��4u��̭�c�&{�������������M�6���7e�h伭��0f�X�ea6`�w�K�A�r��wܯ�I��?��{?+|�g�)7�yq�4�3-3�X�����N��;�S�pZ�>�;�!P�-'����4��� ʝ�����ɐ�I������~[�W}�e�{#N�,w�5
��9��؏OU�-����|�s=���ƶ�/�a���k5x�g��P��U�w��[��ixZ��|$�ڼ��Ώ�b�o_�)��U%���~�$]Ӧ�}}�QL�:���h�z@3����Uo��)v̑�{v����T��&`��J��$h��]�?0�ʋ"�53�O�q'�i���y|�Ӯ(ߔ,!B�.ճ���!L�qV�m��|��Րn���/�x����7��S�,i���Bx[��f��
7�IB����=D1!]_"�}	� ǰ�,��a�����V�)�u�1Q8�\�t�������
��;d��ț�J���$mu�	���a�?&��k�iy��F,=d������2��,D#��~��j���?[���o�vo���Z��no�����A��#����U��5���_��C����A��{�!V�������>m������FzI4��2�D���T@%0-��O�U����j��ֿGm�5a��K��ռ�y%I����"�p�-���־���=S��1I�RN]�ɻ?z���M��'��z��}��ߡ���#��-�a���"��O����v�M�ݥN!Rò0Nك��������"�ez2ck9H*(��׌V�.�����b�Zt��|\~>�[�f"�����(����lF�J�ĖC\;7\�rt�є��+�-��5�T���p >�:��ѱ��v�v(@���E�j��l!��Gp9͋Z����6B ���j��9���X�vv� ���U�݈!��Zn�����Z��)j�Ts�_B��cJ#��	���N�55͍J/�*�<�WF���^2�)s4
L�Bv=�L���{��P�D({\�ln|c�.d�{k�_����fM�%:D��ꍽ3c�6#����ƛ�Akï��Wsj
��8�}���#��A���;w��v雲r�4��"�3(�?�<3�6��-:��d�ӷ�%y��,�sՓ��_:�Y�JJ�@%�(���݌W~�~N-3Gl�W2ݫd����}6�5�����p�1��15��W��?�F
�������<Zl��wsZa���Jw���>ӵ��-����G�~��k�N	�b����p��fs�}�kv�i5�B�PѼ�ey�@��u�E�Rud$��u���o�~��:� IZ�\�0�+�/6���_!:.����GŢ�E��c߲��k�'��@�:�W����qy�z�	&k ˰��J��1d�o8���"�F���fCP_F}�p:Hv����nNk,U����ǫ{�����+J�R����>g-�}K�Ԇ�(U��B�t`_�e-���X�
��m�qS����ey��/�޽���������U�g@�BH��z�n�.:�5��&���	�L��D�fm��qc�ȼw����"�|����?�6��Fy�&r�v=�T��`e Sa(SF8�ٓ�O�OI�v9T?��I⺿����/l���E��j�oaG�R�w�����;�p޲���Z��X٨��P�D�F�h��d�> �ׂkb?�|�I�\@�����p�e��j��Zzq�	ʋ���V�����X��q�ǕP߂:�+�60�5���6�υ��߻w����(����R�<�TQ������%�x��B���:�.�����g�{�
��#[ŰN���{{D�9�Su�J�ʦ'P��X0�J�I��P_����%�|f���Z���{^d�g �
G�3��n��;̜2̗�Cdz�$���Fh�nI���X��+��޳��ڌ�`��db͚J����,x-ʸ��3� n�Nps��-\Q���������B�/j�����s��6�2�2��8єj� ����$		F����+���1�u�S36�0�������J�*��� d�b��$W�m�o�z�a���\�������k�Wl0�>D4Rl%�{����
�����su�A/%�09�������o<��{_S�>ά��XxZ۽ʰ9' B��~!��Uv̓7~$ʤ=�v3��tﺪ���ې�{n���ml"��Q?f%7�2e��8��2���&L�\�Bbq������ԃ��;v�U�9��χ~/��*���|�n�R�(��&��9G�]h{�ySZ;��^�-d�LJL�H���W\*U
`��}l@��yP�3�\X#���a��ۺ{<8�@RM��<����2X�x+�>nN4��:�����#Z@��G�`�f������D#!@�=SgxU8�|����Oq!̢�ۡIQ�<��?=���onW��BĨ�"���ǐ�ߍg@�me�k���|�R�����_�M��S<O?�3l�D#-�H
�2� k6J��	�J;iH���;[��<o�f�{�i���{�)��W�xH!G{��
|���V2.�M��?�BZU���C
�E��$�Lo������l5o_u�oH)�4�V5��iEQ�d�{�����|sC'v����6뾉��]��{dyH���!�����=����
�$�V�����	�B��f�����K�x%վ����y�õ���V�D����;��EM��+�tk/��w{\�y�c.4�!���� ���up3:������SK���Ӳ����L�U����&�9ŀ���|���.L�����D� ��b��#�*��_~krS�L�ď��h��pWo��ۯˌ�ޱW�8yw���㡤`��`��ŭ\�7ݭ���d���&���*m�L� ��8�~+-�����)�c};�X�\?��v{��#;�n"N,�d��(�������kr���#���b�5��I����s><����夫7޽��&l��;����������ZᗺW��9.o��vq������\�R;`[�ǳ���,�{��?��L���秃���D7�T�]�{�(�9Y#X%�蘻{����7F
b�q��j�N!��9�{kþI!j�a'�̶Z�G^k�I�Q��F<���dDMʇ���9>y�(�Ř�ʃ���ա�s��%`����Z��l�4n�pVdP��= [Fg���}@uI�:3���~J�(�M{Y��PQ������R4���v��!���H�~����&���B�D�	>�>�j��)t�Yl클����{U_X$:�:���J�ŗA!����[?Ы:�ъ�� �1e(���Ó&�﫸��L�����d��%�!����ʆrH�����jVmg^�r@�M����%9u���[9|��I ���()��߄�bv�n�-�-G)p=�����n�z������9՞1�3��?� 5��o�RR��ݿu8������ɡ';�[�Ȫ��P�^�����r�jEz6�zT]�XEf��"�.	�wM�q�"���Z�Μ�^���8�WI�8`�5oz��eh�f���ȣ��~� �茽�H�wv�\z�{u��;������\�H|�ЍD�'�Հ��&������D#�{ԑ�s�Յ��QjO�.H_�(��J�+�~�2B�f�V��f���2@Y�\�M�|�]� �O��<S�&�����z!�"a!��7qenG&Z�%���}�Q�ec��kr�Z����x���	.%e>7��^VZ+2N=+A�S��<��fO����/��n<Ei���6*�.����Z����#��o�����sV��b��9�I,���^�Y�l���4������o�|�z�;Q���ng����痶�zZ:��������)��Y�ť��7�\�Fʏ�W?\\	i�6���K�����?U<���?�zF�/�����6�����jh���K�k���i˽�\:m7o�/�_u0.g<"h��.�sv��N��1�N�>�ɒ�U�w�F�dH~�if��[���M���f���7O �=k<[�ZVV!�М��O��U��o�>r���i�C��i�^�[8~:1h��]N�vh��]�?^�>M#�S~2g�B�ZS�S_�������-}}-U�r�j�!��ky������q�&	���8�W���_��y��c���)/�yz5�H�����D�{a���>*�ԗ��=�˘n!�@1z6xCy���wB�۲����N�v����S��:�F����KO����������iyt`?Vi�V�G,�P1D؟�7�*���ZDDI�	�8�}��}ʁu���F��@��߽�O:h*��Вb&�}�&����g�������fq�Z���&}��PEc�9��u���X�v�S����K�$����P
B7�}��[&�_W4�ֽ��a1[���-E��6�����k�M����1��$i�E츺�:@^��e��Fz�7���gAj��|,�vJ��s�̎R��,YY6��&�&��<�l��X*l��*%с���7�����Gs_�V�1�݇�t� 庴ՙ���9�����gꦏ�?{]� OU��rR�PL&�v�aUt�N>��΅��V����}�kw�%7	���7ݟ����N�7�1%���f;��,v'�$q)���S�A�� �zaW��z�?���.��5P@���)Y��MR�������Դ�6�ч�agP�&�[a��6��s�"�լw4���;���oFv�:�$f*��տSZ|����"��vSgX~���޻�}�gJ.�A/Gm>����Q،�ע���>�s�+^^]��s���.���������=�(}@*i��zX��e ��(ў����6��z�G��ХWN��o���8�ZJ/�W�*�>����ç��+��zN�C(��03�.�Uܬ6���m,dϘ<l�Q�����(54q�E{��G}��㋽�����+�^OM�<�����eþ���`����}�N���u���|{�U��`Σ�vv�����x���~o�)0� {�4�g8���b���h(j�VJծ]��ъ�[�U��E�Y{o��3Z{5�&�h�������y�y�q�^�u����u;q��?-���˕u���{�~�GmL��j�r�#�LT�̆��WETF%�Y���.��k-�m�����;<�X�.�ΣlܣGw�s֑�Ə@��������G�8f�Bt�i%ݟ��I3�WxHŝ߱M��v+O���)Y�[�����W���IΑ�sÄ2�u������V��4�K ��h�O��`��i���N]<!�w���Ы@�H7Є�J:,!p$4(w@i#!��Ѕ��(a�RN	Z~���RoyP\���7
)�+����\���1`�$8�6*�2#�Zb:��I���N��i����U{J�l�LLC��@n�e��@�Z|��\�����}�>N���׾�㱐��oV-�����I��ԗ��j�i��a�[l��ۧ894�t]r>�[U|p�y?|w3�r\����=\��"��@ѣ����`�{#��l瀟R���D�-�p୆�Pm��X���s�� ���MP�~����-eC����d�f��*]���1�(���LA�R���$"����a�ED��[���m�.�9��*���$j	ݘaB$�x��']N�������G�;�3\�d��ʞB�L�d�� �(`8�;,6���i��4���½ꅫ!��C���8�oG�%cω`�_Fl0�D�l�1��w@���^�h�nf�p�g�?xߖ�%[SI��a�kBn#�C��>	���t�Q˳���|����ە�P(a���n5��y�� ���S�������1>X˝�BK��ߟ��.�;��'k���L��+�P�^g�(wɟ.��Dw�p���{�!?$��A���\_
������ѡo��9����C_�MZh1�����P.$_�{�>_�c���B�z�ܨ�y|8w'=�y���=�s�m]��;���O���j�FN�|,��!C%�=��r]0cs��O��Z�����4���y2�{i���)�|�'Lq5ے�=*nq(kb*�'�r�0t*^ǝh��|��q��T&T��x���1O��_���&���!��ޗ\Ϝ��Re��9l&�B4����aLUn�à���ɋ2J�QP]l��ٍ=��|x�q�ԛ���x�iP�3B�u,>��tI���	�x�o����h�xvDiOTr���K�*W�P9�fVBiͳ��������s���/�j�Af���4aKi�����#�$�û�?��=��^�A��x�ؠކ�if;v�1sT�P0c|xh�� �3W0c�o�L�d��^ay�Rd}�4��8���#"e,�C�g�h�tjY�3��u��g�+y��좂U�:���R�mqSwq��EME�"���]�3��U-#_l�m�{���j߯ꕛ��*�Č���ZY��������������?��^���_P��x��=�0�x�Fm����eecӹϋ�?�f�8���P�9�54��PbL�ܙ[�ߥ�Kgw��3VnC��w���W��c�E�O�T���7Df뭔�.Ǫ���w�X�*�+7��P����`�vJ2_`8ѩ�
�\5d`e��ueЖ�:�)��]4�灩i��мp�E�"Fk�AOz�-���u��C����N��r��M4�����y��1���,G�2��M9J�N�uaL��Uؽ�j1�즼z؟#p�q�lJj��DC�X��q-oFMU�����KD����#.@�گ���vo�H�N��Om�6�am �̼r�>c#���ULnK�h�y�� ��*e(�-�)��ѧ��GC�'�vU-���v��ѐ�F����i�β�ى���i��//%�^��xF���Ir�n�{K���)t0+F��J9}lJ��N�өE�#Ͷ����v��4�����̹��l�l�y<=���7�^4s�Ur?g�R�1a�n��
�fA��Ǚ���G,��?K�0�Q!�L�7׌W�p�@�]���ٜ����*uU�.}.DvP��/\sc�Y;MD媓��/DV&[��#�j|Q)kL�����}&^v�`�'&��)(�̚�{XD5n���A�D^�X|��$5�>��ޱeg���b-[�@24Q��5��I��P��0��W��6�iR�.���rB��<?�����w�Q'kr��ß�'U��%���}�����J(Ց��v��� �F��Q����{�ܸ���X�M�p��?7��Ʊ/A�p�]�G��� }��̵���?xj��u�����GP�G�"�xgb�y�&�F��H��T���R0��>�y�t�,'�ʝh$+�/�ו�;1�6ހ�Q�v�_�T��&�A'Rf�O�S��º��/�B���%,AS!"��gQD�Ki
�(���L�6˯��S�	���<��L�~�i��5Ã�^>�] z|6�>����*��������P�_V�����B��\�0$+�F�7�E����Gп�/k��"<i�X6U���~�v��F���_x���%֫�%Ճ���e9<��*��h�/�wy�ʮ5��9�>��>�]�@f`�Y����d�n��#��LI|�^4{��?oܪ��sOl�N���h@�.D�����5dS� 6�a�W�8��9~3�gw�Ҏ/v�y+Ag��F��+6�Z:���R�T�F�@��ǡ�D�!�%�X�)2�����̯ɚ��/O�6L�N�>Q�Jj�Ċ��]�6%���t����{�ф�i�5'����+��
�!�f���W�T}��ۦ�%�T��h�����樅הΨ���PEp�.��-�7Q�����j���G�E%3o_�}h�~�g��%�i�t�1u1K�C�V��O�v̡��rN�����j�%����C߹ A*�pf�#����&^����O��X=�?�[t����c:l��y�g>�����=ۘG�.Z'	E���.���N�_'j��We�����L]1�j$�?��>Sֹ8}�#e�..j��?U��{m�;�(��9�k�(,�B��)��U����0/�ZI���@3�xA�qh�D�k�i��js��=T�aP1m��ޮe}X�A�#ׯh�߮�p���9&l�Ֆ�4=[��Ni�Uyo�MV�&'j��N	���z{���i�JE�A�Ճ�,'�p�����q�M䳀}&�roè�?�}�msW�uZ����qm�N�g=�;T�H]��ܙ.Ob���}�����S�q���E,4` v�|�߲��F�����5�Y�g^}܅W�?���QLoԿ��O���E|��"_���9I( �dJ^�ܗ�&�����B�������T,��w/�@H�iÄ͖��P ���E�b��4���Ɩ��<i}#XDܪ�O&� �J.2�Rb�����Q� ���x���c��o~޲�3�� c��6�A�N��J���cI���*T)�{^j��	 ���ǚ�+�1J~�(o��른l$�����`5ꢊ����ʲ��뽣��Z?�q[¤@�\�1�ݵ�^��K��-n���BG<�D�]߾�V_PK7G�r��f�ȍ�q��!�A���ar����k�H�D��/�����>�H����!O��5�Ё�Hz�m����,R=�xSj�Xme�Xޗ�'��K(]���PF�6bg�����H(e}��i�W`=��tm�)��}��R0���6�QW�B��ɸ�ReZ�w�
�a��ycj��A��B�{�%���R�Kݱ;P�5�YE�7�M��F�@�������%�׍&\O�M[�M2�^��)�S�J��%���0�n[,ҔlHy>�^��N��v��1�l#Ω����Ͽ����<�
�Q�X$7�m�2/�Z�v���Th�lr�h��J��8�� &����>�͖�;9����i�m�����Ž��X_�B�v�|�����Z3o���T�Y����Ņq^��pF�����QN2��HuT#�U�ݮW�'��}{v�-�W��J�5����<���^Ɂ�:�y��ǥT��=��
�8�F��K��.����z��B�����up}	s����I~��^1�)��lTx�'��i�U1Rg��Z��sE�\��T�Tq}�%�%H��ļ��� � �G�`<�[�8]^r��P�_�Z1bb�e�/��) ��[����C%3%�|����vmB����ȿ���Ƒ�ͣx�����o�6�'3;k�������Fj7�7C��(�PuD:��輚��}�f�<��ܪ�����=q��nJ�/��R}���¤ٙ��ɋ�n�qY1W��� �Zu��Gǯ�1�O}$?d�'�7��,�]u޴���뤍fK{X���&�=��ݺY��Ո7y�y��e���R���S�0a=�#�A#i�<��_���	A�,�̡��ХR��i�L�0cR2!�< W����
Ii ��x����1.4-��=�����9�,�T�9%�w���I�'u�\E���p�Q<yjY1ߢ�r�����'/�`U��k������b<�)��� �`h�+��B��:�U�f7*qY����?������V�_���%���!LܫG�����J�!�2}� w
�v]���rT����6�I|W)M�o�]����J��J���~2ћ�ݿIL��u�����ћ��%�ʷ���ez���V��>��]ܠ�v�깾�}Li��D�
*�����Ձ���lc%��mX���OG8���MN,]�T2U�M��L�>V�I=�\�銲F#�ո��ל����ve�ʜٻfS���s��iXx|8!�E�%���MŃ����(Z�*��w�´����;���2^EHދ�6�A)��\=t�S�!V�"5� D'��G�d�B�`v����5�r�y>H$�6w�X���T4��F$�	�Ϗ�V'�)	p�ga��L�Q����y)���#T+ǛC5��{sM�
�qW�LMrSd��!B����j[�r��y�g�J&����q�S�n�d5�LX6c�r����l��~�4��ˍ���>���������%d����$�0�q�Q�9�|��+w�{�Y'ȇ����/�x2K�i�(�`?X��߮ő������ T=��b�ɰ�Xs����$1�ş�\�8��{JIs�x�f���"*��0�!��*�QG�9�8���ǼJP ��1�e]Sb$}��nx�K������f��l�l�l�C6H֋Ǐ
�`X��^�2C�750� �Q	�H��`|��qN_��N�h�����4c�ex�-s�k�8���~�dz̕�O3c����O���>WI��ko� �?͠Z�t{sP�� &�0{�RI�i1�-MR�2$�6j>m֒�-i�F[DBݿ���M�g�M	��8$n_���Vy�'b���b<O96={Dx�y�ʍ�vM�����U K��?-�)�X�u�����d�ɣJȘh����O�mUn����;S���t���&zm^�g3߼y�����f�S���y���<v:R���P���Zr��+��3'�帊̸�.K��x�g:ƑM��<q�w�Cs�C�YG��9��Kq��~2X�²�Z����|�|p^g�З� ������"N�q�!�/� R)���#�p�!��H}��*<��9�I鴾U�3V�6���P�ݕ�:H�ŉ�ô���;�c��Y�	4���_�x�a8c�g�&���x!�u��u�βi���!�Nm����V��Â��|P
J��fX.`���Sm{�=�Hy_�.@r!� ���ʜ��׶{Q��R7V��6;L��ħ��s�e���݃S�΂�����F���\��I��^TB�����йoJ���>տ�|x��vL��~�����v��J�EƔ](3J�z���~����&R(竼}�C��E�z��^��(2v���u����T���G���Y��L�{���Kd���!s|�_�/ �|$d�H��>M�
�d-��&�q�
׃s��t?��]��׊/nʮ�ǐ1m��1���#œ��w��k�'m�)��]<�����5@/���\�M�#�A�D����j9*�g�uW�V��Ѻ>8͖�+i�,U9
pS�3�R4٘t�V�6�
l��_�����%Ge�3��Z����B��t:�4�]��ʍ	=�r���~���QZ�k�k�]����Z4n�Om�N��(Y����@�Ѿ�'ぺ�&^y��)=o�'p
�:���$�w��՛ˬ� ̍(ўU�BAӏg�	�|kމ��H�,c��C )T�y�N����\�Cʿ=+������6�55��)t�� _�a N��|D�2Ÿ�8�lnJ����P�s:*~%`JRւ{F-uz���cn������i~��k9V�#���M��B�W���Κ0�њx��;$�J�z�I�����9��=�%����+��bT^���e:�|�����/ISXM�ڒ	��2��d�;O�2��G ߠ�B-3'kuo�!���b�5����r;��`���Q��L]���~����۝�|UQ�Mȵ0��LU�U�f|�mV�W��!}C�D8�[S]���ӄ�%26Kٹ�Fj.s�=����3�y
�����Qσ�w)P��06��M�]����=���WN9aȽ������ꫜl�ؔE2��=i�B�^i[wԔ�y���@y��݊�{k��?^�
�i�Z���K��p�k+�41��=����G�0Sc��A��8�d/>?$2�<�i��|���l8Kni��L�W��Rm��H��qM�^R2b/<W�>Y���F��v#R!)���n ���<�f�x}j ;�b=c�ޚ����8&���"�:}�2U�i92z����y�ԏo�t�~�}���A�%���Šx�94c�"wU��Bl�/�|��f[(��@¼L`�lL���MM(.G��9�����R���:�	��$XR9�zs@&1J�m�)����,��*!	��Rj��9=<0�$:��GM\�.[�Ϲj�^�����͈ȋ:���W�;:ˡ�J�'J�-��X֩ x��r����.��p�C5ͦl7׽�]�w��вDۓBF�2:8����f7:�\�_�sE3����O��R�l��c�[�wuh_������݅���r��K:�uU�7�v�k�N��Ȑ�u+��
Npw�X��������T���^X?���z}��˝J����n
��D�6�ֶ���ҫ�ٞR���h�+R�#�����P�.��~|8��s�j�&�^[�j��7Kr����u}n߂ز�X��p3�x-�6���ul�L�6�x02d�Y&� ��շ��Y~�ѓ"�<�?IA��	S(��#�<�U]l�$�~�↖���;f.��T�m/t�\�ϏR�	M��5R޶��|a�ag�?z�"p=�t� ��$�~��Z�����v�+���ۦ��j�F�O=e���x�BQ\^��g�#�_�z�U>rK���F�"�l2����M���J�v'��+(�ˊ���Ci�A3 ����v�����߼��"���L1�~�׀�È���6�0��'i����uj�ޱ�
���(W��0F5��kds}����Z�1��^�ee2�Z�W�.�u�Sn�e�u������e�N�|�}�u�UZ�|��̀�4���u���RXv�)���ܸ-���#�����%�&+c���R-شL�@g%�&o�M�Aݳ�j�&>���b��
����!yM�'��y�8�P��.�767�!�G���on��e�듭�ڎ����!A,�B�"SA0:BU5��S���qչջ�5.��OYx�3����ٺY��̲�~����#�r�ity'��D7���ׇu3���=��W��<N\�G���Wʩ����/�������|wL�v>W.R���F%�h)~���{L��x�Ζ?2��6$^���t&��yc�!�����������c2���<�5����3\s7ӏ�jR���WO��	� �r�A\Dԛ )<jY/B�.��^����f�����dr1��iC�RB|�$�|����9uR�f����f��L�>/�ysu�x"��|}V) �Q��c�>��v�Z��m}e�ȥ0�@����$`F.�l���o�/OND�<��{������Vx��,4}-P��
&�ȸ��六����]Le0u��`�����}���{�t�Nu  �C뉲�<@R���,*އ��Ԫ��;7������+�n�����x@s���C�\�W�9�)?HX�g�2S�%E����U1��Z��u6��ꋩ�/��P������@�B�V�6�Q��CSJ�7�L���9���"�3�}[��W�8cѷ�>_h`5<���!O˂l��54�9��p�ދJ�3E7�m/�CX���]���ٕ� ��,W$��'V�����@�{��ݠ�o�.����eŪ|���e��l�H�i\�N�]�Ѭ�2r�0��]��Fa�����	ɋI�=�)�3�:ܶ��%�2⪏j�?n���}vs����XY�#�^���O������Up����y��o/�;�I��Д&`����Sl	���|�ӕ$T�Ad�,	��rK=I��C�`ڈ}T$��_�b!]�@��)�T�������%���MXi#b3D�u�i��몎���(�YAi^14��"m7C{9�gq�@j7C���&�å��X��TaK�⚚��>$S��t�[���d,|��f�`��A�toiL �>PEx�8~ȭ'Y�܅��X���j9@ݞ���?�|�'��1���y���F�|�<"s��2V�o�}���-��W��
���E�	�=�d�c�-�K���EA��&H����4��w�9/
�ˍ7Ҥ��Qh���W!�'|C�ή\ʏ�����WF�"�Џ�ƿ]u���T�R2r��`��3q�	�x�M=���;�����6�ZK��X�X˾�Gc%�,g(�LEV���M�����a�0(6Q����K����Y"|�iZ�}�R�|��`��rf��Wn*�v�8)��D�N9^Һ���>&ZV�����?�W������Ց�ZVCҵ�,��f"
�/r���oo�ל��
c��S�k����f�co�c��b��(���4��"�r d�+�P�j8�`(���g�D8�r�BR�Bi��=	���<_Q[Q_,��hF�R��^Sw�+�#�����H@?<e2@2�x�#?�Q��#��l㍪Ƀ�Ɗ�~���6��L�������9��=�7��6H� "��8V�>~�ԝ��Z�r���?�LS�c"��,#����Kl�e'����ؾz�$��\-�r5��I
a՞�|(|�"˓W��w �M�:y8�OT�M�P��o���=�;?�-�::�x]��P֯�YM�9͌�^XC� �F�HEħ��-�M@K��o�)�����u�p���v9Y+��ԓx�b~�E�E�WB7�)��iJo�O������Z3��2�}"�Ld��j��~�=��k�tZy竐���x���eێ;i��I3�~���o��Ia*�·@�R�"�������x:�;O�C�n��]XG(����B���pj3F��=�a>P�^n��p�pF}���4A�� _)�.��S(_D�cyߐ*Q�$�/�W}J�,�a;�����3����%9�Q�y��LXkh�p
���o��|>��]�H������a�������P/���C�Ѹ@մ�޾�8���NG�[O�u�p�k��ĭ�友
�� ���^�x�"k���g�T����R>$�2��|�G=P�h����^=_��ǥ��;�Z�g�q24jS�����:Dһ����!�_-?&+X��V�J�����_Ц����6r� �p=�cL�����y�ǃ�x��Bޱ�o9m�oX�\���3��Qh�,��/��bb�� �
�Ȃ\�Pu���;������Q�p֋L;�"a���*��]�3$�s�rş=��]ځ`끆)�3}gKh[c���[��_��\��N9^_v������?��E�w���Y܋����}<�ϻ߃40~3yO��lꄵ�?��.z�'L�"̯��^�:}��c�	���6"�#& �=X��D�#vR�2�K��Wy�R�J�%�ׇ>T(d7d�(a	
'���(�6H'tm��#�	v�"$�#K;W���X�`N��]n{�a�6��>4G�]k� �O�6@�VRG���$��~���>_�}i��}�B��G'�U�$y:*�'�����~����cņ{�B.��&��*� �m��*uI\�z��,U\�]�]͊���`�}<p©�Pa2�!���y��f�UrM�Pl�!Pw*��%�1'g���������L�ꓠv,Z^�oi|���<z{�n�B�������������#U���*�"�\&y�	�go�P쑌�m�輻 �H��_|�b�*2 v0�'J6��ߠmrB�i�;,!/��g��>]���"�xb�4q�(O�@9��R�4D������.j-Z����%pȉ^�eNd�L��g�T�=�@�F@��κň�b,Ĳ��p� 
�B��b�'��	�����oe�kS-���#{�ZKwN�M����]WT�f�@]dj�#a�5�����ko��wg�@�h��r���ꪝ���	OWJ�v�V���AZ۲x��.��C�t.
�L�S��{����>�ҫ�}�M�i�u%���f��~��O%�߯g�����c=o�7��;���:1� T�ȳ�h�O���1ԣ�7Y�����<�y�=����&oz�(���:����h84`%���ɚP�
�&�D��u�}_�;���c���������+x1��NƞH��D�R<��<7wO�����Ӝw��p9��4WBW��ؐ��W��r�V����>^�.�b	Ơe������k���w\��
�bS�0\�q�ϻ����O��p�b��8ُ����{DiK����H�Wh�ˑ�S<�6��r�q��(>�v����*	Zq��x�.�ɉ���'ӹw�h5�tGp=^e�<�'�Σ��y+����$-���0��~�9=�NdXBЗ��[i��8��8M�E��de�	wO���=��jP�I� �9�����cKS�OT�go��_A�ɓMrs�R��ÞU��9X�=���n-����I���@�Cg��H�4
�����!5 ���j�����=�d��v�˂�>��q����Ai�N�?�o�}�]�/Z�ݞr�B�F�� �Í�-����H��V�����i��'Hd~3h-�����C"��@?(�i:^���=%��Ф�����W���B�I�è����R��KM <�򅢛��#A�P���5�1"}:Hr�{(X����oǠ��~�i�%��9�(��y��'��續�Y�U���ն'R���<W!��3J�_l��j:��c�o��U���v3dO���.���BC;BB��M�~%��^��nlk�=@�d���F��nO�l��.Vaz� ���X��w������b���2v��%b�8}�"p@��}OM;�����Ȑ��w�`��?h�d"p���G-��(r�T ���,��<v'*�h�a�)���s���S9�YPeQ�x���O!�TU(��YmsS���
+�p��H�,p��ȳO�E�[�HM����?�Mmx[�p��9����X���=�Ѷ/j�49�O���w��#���ۓ�:M��������p����)]��^� ��g��z��v�Q�@4����g��2�2�6��Ҋ�\�!��LL����� ^nO+�Pԫ�IG��L˱�kq�ی�������u����I��B/���QV���{����mibX�e�m@��m		���R����|%LP��;E:���K1�{�Hk5q���+���s���r�jbS9xm��=&�m7�����	�S���2�t��"W��d�W� B?B����.8�9����{�����4���J: x�� ��iY{1��F���Rd�@��@�"�T#\�z�)8A!���@�#2~W��aD��������^\p��;Դ��om�@f7�*=�:�&��f��o��m��b�������G�';�z9�p�wBU�U����w�e����Jp�'�޻�g&xR�K{��
#��h��
�����Xvj�*nF���2��%5�g�,�Yd��7Y�G@�' sD�T]ȫ@�AKlՒ�����1��+db��)�X���D`blM ���P�@�`9/���:��(Ǚ"�?����$D��[��As�,�q?6��
�eӯ������n�[��M�{��tE�
�ӝ���?6��u+����x2o��,@P��p��=�͞gm>��:i"�z2�aU�x�"dT�=�a��e��Ř�*�z�SC�Z�N˭.�� �91����ZuЄ�'%��/�q@��+�ĵH,LH]���wK[`����ͯMh��P�é�g6:�3V��,�M�MN}�	I�A�w`�m.�l�1
0`e������'�� M�A�+��oU?/>�i�ND8�<����Vq��Jr۫i#�����L�1r���������//��<Ï��zU���n�{�nm<�K��"5ؽ���Q�U�9�5E��N���JUt����.5��p����a����@��hN�5�ˮ���b�R�����R 	k�7O��,,w	�t|TA?L��RxM֔�Z��_o9/���'�U��ϴ���`��L�vH5��m0$��zr��e*n��H�(\k�˽l��0��i9�7dLf؎�M=�dK�S��X4f��� ��P�qye����vH���S��4oD��}�~�ѓ�d�3?O( R�(��p���?��mۡ���DlZ|���3��A��S��O�3c##�0�.C���2�H�,ajps׷UϿ=�w�	�c��hжzr/Vh�2�<������B��yA�#�=Z�ö5�y���rT��9�X�m���Ϗ�n�q�uH�᠔FW��Ϳv���AR���pz������ɒ:�' ��EGIh6��`��gvؤ�������=�>��=,�q��o��O2E�D���(�w���G��a]J9�?�J*iL��j,,m�u(U��`k�A?G��'�s�Ӵ�+^�'�<�-ݨ1RORwR_/~�T�z�����)k�-K5��-� ��
�
�a���Y�V�%��v��A)FU�<R�u1�j��)ȨG�&de�48%��iU����>N��j:����HY"j�ѽ�S��p���oq �Dq�Q*��6��liW���Y����/�����������-����m�u�.��/?tD��[��4<��vv�e���gu?=� ����L��W��O�į�Y�"����8�W��;,�%�+ޟ7ܽ�u3�L�0������)r!�¸���5���Q�����W�26���w�S�����i�`�)n�!��|W�T����9���s��u��e"�P����"�����=�1ƀ�"9� �g؄�1	��}��꾟�/F])[���PE7�C �f��tI�AM�����)\ӝi�R�lV�ӝm�;��zSQQyok����.����d��S��N�W��S5��?E��5������Pp��B��O�PZ�-�}p���o[D�|�݇���c�8ri>�@�d�.5��������i�h~�dy���i+���S�2���� Oj��g�%�A�l����[V� M;��h�e�J߅�wʀ���/�ŇZ�|]�q� � �_�=��۩��)ؔ�<�B���¸��
���u%�����F�o9���blˏ�XyA48�$�mִ-��(��ioL��MT�G�,��~/��UX����Xt��f-��H����[#�K1|'���	JU/r{'�o��m� ��#""4��e��s_�޾=�����Υ�|A#1�B���82��W�.��~��~���m� �T9�� E'��9����*8�$x��U�{���Ҵ�L@��Rʼ&U�T��K��֑��	38�[��"7o���Q߿������`S��TJ]���c�d~����o���F&K\6��.`U���]7���"-��N�D����!�$`=�Lw���de*��ݦ}sW��f��7-eV��?�8�o�8�?!^�����H�L�[U[������s��r��z��8r����N~�@Z�e����Z�)�X�?hoV!{Q���HN|>�詖W8�W@ 9���К�l�QR�'Mr>%����\D��#$�����3�b}���s��~�_�!�<�Τz����������âɃ.m�p��<�;XZa���.��X�Jh4�u���l��9(���Y�;*��b(Я#<������${�4�>k�I�X�>�~��):��9r,�ɇ[s}]�wTo8޾~�t۠��m���s�K��]*�Eۙ
ӷ#9�_�(���������#�B��M�_�M�}M�IK
��r��*UN�7��*yOZ����#�cr��6H�dp6C�*)&s��f�?�u� �){���A���m��q���Z{{�)?� ySJ1m�O�6�Ȼ0���e��i���Ln7��k;��J���-��yA,^�-L8��1\p��N��$ȭ 	���[J�
�y|���iL\�0��l-��;�p�L\}�|S'Ȅ�z[�~6W��i��N�^d(_��_|�oq������\���a����&sF�Ph�j
�fN|s�l��r�,U�U���<��L�N���L�n�M���Y%JH+�s��½q����V��_+���X��ƫp==�6y�c��,jt�TA%~M���Pr/̃n�m~�u����B3�N�A������o�h&n�8}y��r����O���?#��ww{��3�r�v��_�}����H]�� b��<�8.��nԥ4�'�������D���չ�E����_���~|�m�t�
O������]|��{����j�9��]�6��� ��(�T{n ��AD�{�R4Z:�����9־��;j��-�9��&�7�����0���%EKS��DT���wJ����c��9�N�_����§3�l�ۈ�����J۹lL������(�����4�-��Q�#�#u�����#t{��"����������_�m��r�eO��"���?��Ö���o�vQC���)Z6**���@fZ��ܷ�֓@(K^�c�3�u��H8KP�z�X
�JL���&W�4Q�R�1��{��x ����m]�ێ�`�n�0���I�N��ꨅ�ۮ�2(lg���~(&�	�Is�F���";U��;V����Y_چ�I���ۘ.�u��ݛ�/�j����4������2{#Y���A��/'�)>�~�Nҿ+��D�|��W���r��Ո�k\�%��i��n+~�A�ġx�HQ�,18�:%H�A
 ���eq0~/3�p���gB�6R��fMv5ݺI�аi"���(2��@����h����9ʣcT��Z�R����⥩�yez��w�ő�u��Ɨk%�>�ʧ`j���VdAx��ji|����Uc�~K[�� ���
���Ɯ�$�$��.׫��_-_�L���h�����|b-��y������Ҷ���[��a�8SsL����rH�7g�� ֭.g"=Y�-k�uJCX�*B��� ����St��`d�vݦ�utp���LV^��|��U�G�2,0�﷬/�l����jLlH%^� �͞��T[��طL^x���l&�Kи��q��R��dt�hׁ��}�]� ^�Ҿ�����޽�:�7�w�+�؆:����̌|��D�������R%�{f5����X2���PJl��  ��C�,�,N�<�d�
�I��~C3>yԕ���]@V!�dm�@x�Z�t^'l�7��
d��tl���}�9�q ���&PU�lV'4&�g�`��K�^t"�/�'�_�E1���-�d�}��hw�PȤ��S� ������4��c�iq	/M}B'���9�a��Tb|w�bC�]�)ZoL�m�������yi*?���n�i��o���+{a¬5��6���i��B8�k1�I�'��F^a�LS�q���!m�[)8�wYk{�AJD�J�Lm�+�pmL���X������Z�5O�������rq㰦��ܛ�7��#���cGr�f0)�R����(���_��7[}L���^�vq��nm�����?^�}d��>W�%�܌���O�j��V�	�<��H8&p��w�ۏg�<ZU]O7��vE��x�KI�PwFjj�g>j�Q�?�C�x+�6�瞪�b��Pp�vhY�w��K��W]��
�%�������M���w퇂��a�[a	��b~Zz��۝�A	�珇'��Ŗ��jl{��z0v�SNB��^].�2J�-��{�8�;T���B��Т;�m�풷����M�>��᷻-�fc�
orP=����R�j��Ŷ�����?C��+���y�v�Q� �U��O�M�rAhǐEQ9�",&�Д<Q���E䧥��K �/�F���0qK���c�p[�Ƭ�w�E�Oioe�G�2C7���4H	*J!ҝ�t!��t�� C]R�ҍt7��w���9�{�=��5�u_�������*�j�ƌazCz��}����J"^.ҿ@-�뙋�GM[�6�H�osۛ6��9����"jf,1r8����ƅ够%�ܒ�7��`ď_��Bp�嶤�n�d�&�r���$a���O�n�_���3~]6���xfQyCȓ���<���x�X��)�0��]d���y���9����bcbNb����Ƿ�����4�[�9,�ъl�u�+f��
T���bM� ���:N��~�y�f �J����YCCC%g�}�/���\j�5�}MH�b�>�ί���ը�+*^��9)&4��
B�-���O���]4@�G�O݇$8�D�9@�BD_^_|������y:��gѷ\��տ �ՙ�|?�x��dcc���lA�$񲤇�#�7���a�Y_Rq$s�g�)��ڴ�F�d80Jyx 

�M�`�5����<���L��Q��:�{�LkAdH�d�Ŏ�}^�u|�\�r��d�������$�Uɰ�{���(%��a���o߱)�֑�R�oYM��0�C��kќw�(�6�~X�Y��v�Q��ӕ�N,�v��צw��H"w�K�6}�r���b4Û�`+��\Yb��;�>s�>������[�=��ڤ�(Y��� �b� ���Y���N�5�����v�Ւ
ė�_h0�S�<�19�К0Od:�� Rψ{���q��,�S�;��Jg���%(Խ�L���nu�Xg@dڴ;Li	5� ���'r���V�%{]m�O��T9�G%�A�5�@ahB���Wi�C�n�(�7��'�W�����k!�}�kyoC�wEQt��� ���)u?\���d�T�x,���`m�@���$A2|4����{��M�jO����?Hȕ�%�031�:���+��N��`h�v]}�_"�!H���1> �hR��������/v���~'K;��:U��=�J��[�fOs�;�Q�GL�!���۫@�Y���NDŗ����I����̪�Q�r&�x,N��V;[���|�Hx�}{>u�Tߊ��=&sQ��;����H���z5�+<b�Q��5b��-Wd]��=����O����?`O�^�a� �/�^�E���RGj0�%��\�z���d���<�����:����3p=v{
A}�:83"�v�O
�G�ϛ�jp���e�᫙a����%��7@?�8�~�w������3�������Kg�p�d�p�n{��.L\)Up�F��*�a5Rx��	�+�^���׼#��i�Q꯷� W�k���Z�:�JאF�‽ɑ�#�kd��:6���ҹi+�:8e0�zO�t�e-���1�P�^�OnL�w��k��#���.��۵p�rh��F���.�a�+����芘b�`:8�d�Ϣ�ԭ,��O�U����$��-��4����N�%}���0��u����Ռ�B�e�n7��w�%�ٓ���ii�7w�w��%��e32�j4���T<��k�`�7EkA��JW�I�:&~}bs�D�O`�1���'�����*,��>`�G)Q�]Զ�d��W�Ts\fuj`[T��(�`���9�c镇��ԑ���3P�ǀ-[%�e����&9����|Z�1�1/Fr��jذ�&p��t ���Jr@2� ��y�@z5� ����v ������t�eVx���q�X�N��Q��,�1�i��n&�C�3/g���Þ7��Y�J�����z'o��0p�o0�6��J���D=?8�b�H�w�� `{��1�vk�@\|6��r�f��tHrQ�LG0l��l�DX���HB@��L��i\��YW��&�����	y.3�D�u{s\ޏ��d8	�z^���e�j�a�\b����"��N`�w�ϧSzLuW��O�� g��w
�--�&�l�6ʙ�M��5U�5���c]�(��m������%Cb����+'i�6Y�-��m��l�+����$� x+��_�ͺ©��~�����<��:0<{q�"R�n�����<���nc8���x���r���0*K�NE���K;&f6�}�`�t[ۊu� ���MNR��7!�:���]~��`�����GN��X���:W~v!sIȓ��v���P�)��U�Y=�:�|�x��WH�
�p�ҚD��������bHh���U�\���k
��7�C�}�ú{�v��BnOD<��0�F�� l�3W�a��  fn�{���"�.�j9�?%�e!D��� ���B��l�(ZE>Ha&R���T����H �ͳ����Vl.86�W���v���6�q=f�7J�vR�G/ �Y�j��@�H��M��0h�H��DG�A�SL8�L�?5N��R�)Zm.��Q\=(~���6��I6 "��E�����2`d��)A�������!�%N=�>,�f� ��n;����~��ҏ	���w�k_��4��vb�7�~\�`4�ޞ;��]�YO�O��]e$��׍��h�n(�eZ�k�Ѳ�s[p�FN��M,xn�Lh��n(�L���l�&8���p-�A\�v�_��)���C���҃Q�6r��E X6C~n�Ǔ0  ��Mɍ|&I��h_���5#���[��Ȓ� �5H��G3���,�e+"Ȥ�GHyyOV{��b�<c5�2����@�äQT%#E�6�����·�O�ah�6�~�i�<��m?rW���l��J���#���1��
����U8k�i����P"�u���u�H-��ǛVtb}�j��Z��~�v�?�h9'���z��1��g+;k�S?��gf�z�	 ����\âf����U��~<�K��:�׬kO��ZO�l���y�Ϯt�D�w.Z�0ύ<��͍䤫�"�������e��f̈[E���lǔ�d���$;�^`��2+�m�6%	S�[[q9�}%��#�G�t�B��h�#��Ѵ*B�]Vt�wph[x^h�&?�}������U��Y�>�=���N�0y�������؇T��"d���`�02?�p�����k�e��o��V#�g�+�nlJ��]`����Fx��;�62(I{Q��sV3�:�i�����!c�0��_S�x���wA�-�wLߛn��Jd��K��M��U8�aB�S_�2��IbHWc���Y�ylKXM}�`Zf�_��0­�I�+��W 	��b��G{ti"��X���_+�(��{��1j^x�M�*�+_�Oo�ſ�J��a�e�e�����6��<Jfɦ'��{ �7�`�׺�WI۔��#�a�F*�s��xm��[$b���X�[��L(m�ʲy���\[lηV�=O[�ޝ勻,@A�"�;Sȕ�[�%���<���?�$͕�� ;�����qQ�YiEmA�P�������G�^B�n�w=�R�ɸ����%x8qK�1jSʵOp�� "1���q�՞-]ӄ/C[��+⑵���<J�-����g�d{F~ߨ\0�"�f/Θ}@��'�̮}���FҘ,뫩[>���n�S�si��FtfD��_%,�mb�ß��;9�d������8�����0���yf�JB�h�ޅiΤG��@,����L�j���|W6���f,���_�����K>��܄��F�kz�]�fާ5I$�W>�p
�kr�%�Ӗ��]�X�g}���lK��.�����\��F�RTV��4�"�;Ԭ��^Z]��$,P���t`��-���D���M7��	d3�I��o"u� �1�g���U_}L{�`$g�t ������F`�;��/2ޓ��g.������C_�ʣ �q�/}�Q��Uzy~�������L�x���*��#��D�����AW<����32�y�"�-����$^��uB�!u���:n�5k{z�/h�D>] Lڕ+��΀F�%�������H2��1�FK���\_r�f��4�H�����f�N`�i��n�ot�j��z+A- �55�#
�G�7Θ��\�JW�D/W޹k��8����蔛.e#�N�ϴ��vc�mΡ%Tf"q@�{�����We9z�����*�d2$����)vZc0Vn��E�vg� Ԣ��l�9������k�0sbc�&�
iQ��I�ʔ�'��Ô���;���FG�� Ɩ�ԃy'B�y��MǤ���J�/#�Ӡ;ٖ6��fְ䅼DÝ'~�0��1ǩ�-!�OtP����݆]���{Gf��F��Z���;/��_q7��k9_�[:.-�v�Ř ���<lB*�<ݠuG�r��,&��i�쪴��p�����}i��,أ8	�F"��n�p'������������4�@.�Q��C�-7'�Q����_���-@�y|-��dΌ�@Oȹv��ǺU��[�U��NԎ)r7�w�}�J{�<��t>��9ia �o����mY2<����
=�Wm����Ck$\i���������Y9Z�o<t�;Z��M;]�5�f�Ͼ� \�a�>	��lkX�>e%��=y�3��K�o!��]2ޘKÖ?oV���3�[:+�N좤��{#��ź���J��*L��ݜk Y���f�	�z1�_�+�2t�=D;�|P�,g7gQ2��P�]:h
����	4ML�9.��X��:�n�6j�!�-�����L|M`|n1vqA+�37�f��Z�M�0�0I����z���W��ȭ����7_t��ά����a莕��Ӹ,=��E�I�� E�cj�Nc,� �pYҖ=�N��3�6;HU���]�f��"'k�{>!ˬ���+�w�����:�'��9���]�}~J� n�uD����� b�WNa���FGgZ�S7�{GX;��Q^���p�$�+��e���1�$�򓐨ө�6�A[LU1�KD���=�س����'mElc�pN�nH�R�r�~~3���o&�p���B�z腪b ��u�e�����p^|��軥*R����_Z,x1+t���)����!K�64{_�VcQY��p*x�F@��l�2ڐ(�Gǌ�e�5���V��;������'��Λb| ���K���>l"v�����,Tx͖�vrAe�6ڳ�!K�[5��嶢d��ic�f
���Mg�~�ୂ\	\D�_ڠ���NT��?+�d�3D��S,���z|G�B�g�9�S���6����k浘Y�~?a��A��??�B�I�w������T��zg���q*��XX_�M��Vc�ԚZ�`S��z��aؾ�y,υ����I.q�2��\�����F��V�����ϲ����x������y�nJH��g֖'f���2��;�gc$�>sk�p���O�"�_�д̋�����4]�6�y����9�Em�Gɩ�;��!������A:���f�$('t~�N�V]jc�b�9p]�r-k<2���ޛ��(֫��+Yѽ>�6��Oul`�[ ɪ8�h��E0���������'p�����;xF�Y��O�X�*x#�\�qƒ���z_�����/�Hk�t��t����ղ?zdmf7j?A��mǣ���=��E�^H #��k���k*q	�?@�S�����ɤ6/Vˡ+cQ/��B�G�����qO���h�Ũ�&��C9x������?���(�yS���WM���Α&^�ֳMi֋�֟*��>�}h��aq��1�&�;Zyb!����M��Rq�ij����� �"��uδ!V�z�A�IU\/�����������ҁ.S-r�Su�u����ˇ��T���.�]7�~w`Ӻ���p���f`Q�ۉ�?�/a?�[&Te���_=�p:$�-�| ������u�U�K�T����0��4�¶�rc7��#�5KU����'��5�@���{�
��gb�{�}6�mIF�;�f{�f��|N�Ճ�s�
(7S�BBh	7�5vD̮�b8�m�o�/���z�SF��V �$Z�2Aţ��uVo���8>sa���#��J�|�ܥ������>�ڑթ�#�ԋ���~�էSB~�La�Q���eL��E5�Ϩ��[����D�����J�'sF������=�`��s{���Y׷���m[����n�&�V��J,U���w�ݦ+�s�ra����E����R	kd�d��n3|��>^�]T�5��]���p5��s=�����P�|���]��A��)��FB��|h���Z�� "W��Q��1��2$f�٠��\���"b��
�^���i���0s��� ���rQ��z�.�ri�|��bָ5�ޘ�1��0O�|p10��>_����B�
:$dZވ��Ż'zf$�	�5�o�fz=1C�`7'G��q
�����Ι��[�_�(����t�J?fVpA)�����o�m�޾�4���W�1�n�ІFn��*tK��n���������B9� ��J�H^golN#��G���F�N"�PAX﻿./��Qw�`}�jxӛ�I3+�L��5-�?�L&Z\����J��I�2EZz_�䢙pk<j"SflK}(%����|i��z���i����3���TS�?�$S�3Qg��=x� �e�U��_k�Z��S����MX	�bZ՞�����_�Y�\i��7��_���o�Y�\�X���0PI��O�:�'�3��X[�Yq�fmH���/[X�	�Jsssw▆���ywBc��1�%�$鳍Y�]4*oДWtU	j�F���gF�
z��Z��]g�x��F}6����p��TH�ue'�_K7M��&#Q��a��.���d�Ԛ�,}M]��m� wz����Ə�u��ӫ���Ϡ*��%�=���RT�Z����న�+#���1}��]m�#��`ӗ���W����L���!�=#�
����/��r�.bIWpQn� +HKMMM6Ff��@]0��9��γ��Î��Q#Q�^WlV��(�)B��I
���ޖj=k�r>J��C݆%i~����A(8�ǍFّ3��e�P�	+$�x0-	Ɵ�&qz`���� >az��EW7���r�_56�V�7/�}@-�v�ޝK���8M�Eо�)V��Ry���vn$g@��#Ε�'ͣGM��%)%)�p�3GcL%!�Xz@��Ii�Ksm�
���4:�$�ߐ=ԙ�S�	��C����9�̮�9-S�-�M}��%/����+�>+������G	�Fd��>{<�H�F�ͣ����
`�����Uֱԏ����OL���[�Sn6�Գ�cEMG�{E����Ê5��8��8�Ҹ�����5?�E�Α��ԈL�L����Iu� ^�1'F	��|9A�#|�ؘY8"=EO��lw��TwW�=�2R+��&�&cU���
���l��
���;[����O��6���n����.�:1�*G�u��������D���+�� C�A�RM���
��} G_�?{S;��BA���<&FA��&�4a��B�H[WO�)#�
 z��rM�v2��1ϪI�`�$㉵��%{?���9�ԏSl���wu��/�I˷��3�����'l��01��P�'v���G���<�u��6_VF0-�d+>��mN�7�����/,�:ݥ�P��u�(�b���"�z��N��*�������Gb:Lu

�r�B�٢���IP�y�Ϊ�����@Q��0>VL#p��e+~_��6\{m��U�0��'�	e:��*x��'Y��/퉍����i\Rq(a��� ����,:<�1١�$���BV##�Fg�T��8�Y �[U.�qUb2�s��w��o��$�$~���M��E���c������^&*	��~h���;�~`0!��ᬤh�?|��+��k4�D�>���$�$ꪥ���L�k���7�_�M3�B�֠��������Y%5 �Tp��8R9�ʚ��K+��b�����ۀN�7������1��0}vI����`��:7�5�2�.����wO#/����k��Dc�#ޣ	��v)��~��~�W<L�6�F�v�����bަV#�λ��$�_5犯��m�c[#C�϶�I�;���ng���qqep%psAlǅ~
�9]I�U,����y�x�I�?��������q
����:��<�R{�FJ�+��$蜱�S�����_3�b]~f��G�foR�|��Vî�Q�?ejU >����Z2��RJ��\�,������<���Fwf���%���H�F�ܷ�6&e/;�+Ρ|+��"&ܺ�F]�d�C+�V�$�ڗ(�����tQ��^�,�����ЙL ����]Q�E�ĨaZg����R̒�
��������V�Z�)a�J��7螉�T=��$rg�j']����R��~���'fh�0B��5�eٴ&�?^����kdF���f�h�� ^tU�$8�,v�f�B�*Us��"ގt|}z�HR�5llWc
*-�QM<�����2��Y���cm��'���YZ�ܙ1���CC?,��76�K��p/؇�n�oC�M/�PV�4������^�힤s��G}:C��1�}-������G$1��
hMZ���U�}U�F����� {VV5`���c-<Wk9�~�B׹S�u4#EN���� �$��?�k���+R]��C	�.����24��*�=?hFK�a��MnR���悌��o�B����`��O0N|/�ތ����N�	�I?D�>[r��a���]�ͪНF���y�Ĥ�2	/*r�eQq����[�lY�nXp_E�T���Y��?G�lʚ.>�=�PJ�� ^�:繙�p1�!���
gç@��8	 n���jK��c�=5s��(�[�b�i�%b%~��$�4�$�_����O��u�?_ɉ���Yd�jl�� ��O�����1���9W�r�Z
��E��y��0��Q��)�F����/�ȱ��\i�A�$e�F0�_xGe��*^P�q�|�?��6<R�ς%z��n��
]�N,³�Y��l�D-|&UvbIwQ�)�.��H9��z�F5�zpR���|�̻Ɨ��w�F~�~k=��k��.��}j۞h���� ��)#��@t2!�ڀ[���u�U��$���A�]���4ge,CO��W$�bAt}�{!Jˋ�@v��B����~	��p��#���ł
N�ŗ�\����"v��;�E��i����zʰ�������p4g�za��3��+�g���S7��d��N��{������|}��զN�
�_��-kYLB`G�q'�4vԴ���~����F O��ޢ;#�¿�rW9�,lờ/~[(�ZkZ��sw?��lp\h�g��x�^�q����߲8Ez�2q�Z��!6&f���u��g��%rkl֏j�1�R�M��I�������0�̃/D�;�;O$��I����uV�ߞ��(�,�Wfz��dn'Al'�9P���_��SK�(�Z�55�/�K�r�=����*��(\�%�(,-:5�^���KX*�I�~�O�����Ύ�tT���(>$1����4�6������V)�7�7a0��<|�/�.��	��4{��w7�(OǕ�o����%������~+rN:��Ꮨ��2�c$������d���~}�Rl��n+��vy�?Oܧ��2<�S7^�T<r�������uL�	���p�"��;ϯ�c���f���?@��=k�ݟ��t�e��.�Ӿw�kI�J�IY�y��T��U+��$A�ٕ��n+�}Q�o(��3f>�N�e�<IQ�*L�u^C�=]6o����5ߴ
����1���^w���}1��v�4��!2��2��GY:_���`
�-Ǻ?X�� bK]�I��ǯ?5���Rp�TH��Ovf��L�ܕ�(i�-H�}�tq�k��3k�����?��3�1,S�.Sru���~8��F�|,s����NK*����9��qie����ܒe�垜�S��x��u{��fާ[4`�?KH��r�3J�7}�Ys/.3]��d�ɾ�'�~�������랐gJ�l����׬�:�S�ڴ�����K��61\��p5�A�Ok�(;�U�h%�����!'+4;f�8DHH���:mݖɿ����sy��d�ЇşL�0���A��s�v^�n1tΡ�z�k�{�9�N����jJW+�T�>Y�N����e�L�lj/��*u,
�vC+4�r�1��-�[;�,�z��<7��(#]����_.����F���c�.�Z�C�\$s'E
,�^�~S�(M$hm@9=��V>��1���|7v�븓� ���-r)�)�^Tڗ����T�ϟ��bǚt�96�m/+kXVI�-D�s.����}�<�B2[���p3�[�=x�W�~C�f�@c6-Ц��	jw�J�\��8B��
�O���FFp@�R�lFϰ�+��/f,�G��@Pc1-ba���|	Yz�kP��3�e��3��;���M{�,���?=O+�o��k2�)-��VB9*���GA�A\�B��� nPشm"?X�]�;fV��\��ҧ"&+��S㰞����{�l�?�]f��wPR���	i(�%8(�3y���m�$P^Zzp?#�b	�UY�����sӄ�����Ph���]������6u�\�����&��s��ӉE���M���M/���(>�u{�^����4�"H�ۜ�3������}D�o���+��,s[>^��4W�u ��#�ɲ*�Y"���b��Y~w9�l���6�>�|�	�#���̲���߭O�76{JBJ������+y�_�|��5��s�J͒��TN-!��)����_gcߙao�Q�X/�7��E�&�9���+iEfJ���MH��,�m�����Y"a����%g�'�fW.*"L^aG�&�p�B���5;�>P��` ��Qa���WT�b�8�H���m�v� �׫ z9G�W=��?������C9D8.��<�6_\�W�	���<'����!I~f���-��gVc���L
@�`��׼m�f���&����"�"l�ݦv�C*�o�{&�<&3D��;���.M��w;?�����:n[���%7 �ص�Q82�v��ċ��������j�˹nM��F��h�[\�!	��hc�=�r����@��BmI���+����Jk���r@���
����W]`�e����5��7X�\��`.�"��5Aϵ��j��J��F�t ����Ғuہ/�^{�F0W6�4����#�&�"��e�=���@0���y�%}x8E�K]������|����E��?>��n9���P[�=������>�7�vI&k��8��a�N=�b[�6�.Rh�@�p����i9��/�0���ϼ`z4ƞu���D����X\�ET6��=V���/M�P�n>uV��0���e�O�u�ad����������!��*[|Mf*,��u\l�n�s�	; ]��0�>�O�zE���4����va5J<C���I��-�4��a1D� Ů+��$�-5�Sg�W��Q�v��G�_w.��J��]�:�-�%�b��)�5]b��e;T=������N�z��O���{�,�����Q���`��>���
�^��rϰ������k�ar��U�sZ��I�;�u^r�+�;ɐ���cW�����t*���D�o9�U��e����{}�����4�: ���G���
Le�Y������D�x�Z⟑�1W�9��*��yTa��v(�����=L��Z�}���#D�D�S�ʢ�f��ʌ�L���*�96M��
��M_��8j����a_Rl�͛O����=Z[sF��Y�As_�۹:^�- ��7�O3��ء3�:�U3�Z�\%�_��vW���H/�ѧN���u*���B�
PC�q۟1����x�:"SqF.�s�qo�ܱ���i����j��a/�1ؤ��oqn��i_2а�}G�h�������.��3%�&1-���Y�	��)A�=��K�OK>����H{����S�?���r:�OŎ�_ ��ϲ?���f��@߀q̓���)��&�P��t5�<��U� qِY��ސ*��)!�/�fg�F��Q��3��j:�X�Ёv/0I$���Jjwl����ߡ2+�֙Rr��3a�ow�5JǇ�
c�>rF��9�	�Q�H�X�˶��^o�l{���r϶'���U�=�ei�p��S�7�b��x��_/��)g(�����pfh�� ĭy�ZvkV�
��3uc�dKB�@��!���V;*OD�-$t�-�P��仯�,3	�8Xş�b0�k�:J(�y�Va��;Z%Q��������J�B��|W-������RfK�^���t�K}a�6���w�]b�h�! �^}4E�'�ܗb��Lu���*����L�ӌ��<e|c���ȼ�g������w�Xlfx;֐>���_¡�k�klS�+��:y��L���V���n:�s֗=���U������#��W؛+iit����X"�����7�-�չ����^YםQ��'`�dȶ�y��2�b�/�!�e�Pb�ן�ސ2C꜇�^#uu�,��1�lS���F������f����wy��X�$e��������_Ei�M-�؍�,9�b�s�U��%О����V��J\�{f����1o��ˋ  ld ��2+�U��P?]���ac���$+h �q�������,��"ڋĞ�n�}1c��?,�z*|׵�1L:v���&���!��Q�cjG�?m`���!oȠ�)NF�՟d���V���_䁢��c��(�j�^������84��~�v���������^����.|})� L��(J��B�޴2B޳ ;�$���z�<S,��`����f*Y�Z!|u��f"�61�C��E�1����Y>��3 �+󑤘g�m��o�;��30Aӎ��X�3�]4/{[cV����c	���X���zK�_����>Y�g)ѫ��	P9[�Ϯ�I�!-�?럸-�������d<��B2�-A��<���ZЏ677ǂ���t�[�1o���l:���+厹�x�rA��3:LK9� K�ޯ{�/A��Wg��C���� C7�҈��iњw�)�/oG�.w~�#N�[��෈,_ߠȨ�a��I����V6�����4�&�E��y��������o���.a���]94���h�ӿ����۽G��r���6E>���oK���PK   $xXN�v4	� m� /   images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.png�{eT]�����ˠ��Kp	 �Cpw$�%H ��'��Kpwܝ�y��_{���9s���vUݺ%OU߉��*��F�  0d4  j  � ��B:��Bt�R��`�H�oT=w �P����S�^�����t���6s�X�Y�Z�[8;�譅�(ʼ��u�����.q6�n5&��h��H��tҠ��_���o_���ݰj�9�j`@LT_�Z��d���BX��%����T�^�O?�ڻ������;�^�t��#{{Thm�+��j���J;�?��G,d���)���'eH8����%cG��q,%5'��O�N-J��dj, 4��v8?Y#�0Ӎ��?�`.�V��z1�O�������{W�8�^����ap4/~b^���P��^���}��@��-:P��:{1��ΑW LQQ���Z?���U>�Z���N�1C�]ɅS7�HM�3���?�Y0��sZ�ۅ'� ���%,҄nl!���wD���`G�b+��O�~������)����,�J��z Rɻ$�-�TR�*Q8=g��?�Ѵ�Y iEH$#'Iz�oY����+�a8=��b0ҟ�B�T��}��;5ʻ�;$"�;W�P��$⛩�4�_g�,�� (7?�Ɣx0@b��awr��`��1hdb�Ծr����Cq�Ӿή*�Ä�݋�q����LR��\�v�Bo�`�z�̐��I,���F�4�!�����!�
@�p3O�ij���0.����ZeE"�X�%<|)�ؤ!�`3�2����a�ƈH?��¸�$�� ؈�H�QGjC�T�ژ�B�`̄y�#����vm&��"��[B��IL����g"����RhY-��C	�
�I�H�VAt2�w
�Z5����얜����e���!V�?���>4���>*$��H՚�n�	�RBx3N�K�#�u��_�u�a$����8�d D��1�J3 7I�*E�ưdB�������ʠ�DJ�~7�S���yj�d,�8#V��K����������,�cʪ�c��C�������b��Z�8]| d���f���g���sj�=�� ��x��!�&1�r�Ӕ�`�co����#��&�Q2G	��~��^klQ�0>�s�5d g�B=�d�H?�JsVP���/�ama��&��?X5]�(b�Y���ӣ@��w���'�.�7igi੅�)0��VK��E�i*W]�Tu;=�,����?��7q.N�;�.��ڴ�[P�B�6��[T����*.E��ہ-��'_sI4�Ҡ����:���=8R���	*�+��t�}�k���7b����{��>҉"�T>CG����WV�Z�����Qʈ��^�	�?��9�̫P/H�"��w�Z�S�;WT�x�6��:��I�R��E���� W�}�}�{�*К�ì{6\m��%k5'u�A�lK������l�	u��4�x�J�r��
e"
��ו�+)�3�+�֔�OhԠЏǻ��qF
.�^�TȦ<�dJj�_y�8=r�v��g�E���0�ۆSkJY���{��u_�#��H
߾��92��8���� R�b~�4u1p�iF����".pP��j���{�<���ٿ��Pu��,���t�ڰ)կ����ݵ̷��xv�լ)���;f��h�N�y��?���=E,��&&���;�"j2y�0R�H���)d�����m ؉����3�.� �U���ցm�l'�2y�1����&T�70vႝU_�X*�X��ˁܟ룽�����<׋y(a�Bᇇ��|�է�/�Vē�'�)�o��@i�_Gx�����I�UeO�Tl��	j��#��Q�TӃkw���G�C�#�X�ƛ9����2 j����J�xQ�eC� H�X�f����t��tPԯw�A�n�r�7}���R��uNOǈŜ.�{����U��	��z��잤�a;��ب	��2;�<�U���[�0�6CZ�zP ��$�;�k���1�����-��&}��ܢ�}2Bsh�쫠R㥭=�?��65$꧲
�Ɏ"|��b��{����|���M��^�$�0 q�$"��Yo�Mp�+�ڊ2�#⫩�+�>�����J��t+��)�W<!��K<^�>�ې���YO=����Q�%�rpb�Q\G�vË}il�
;͕`N����Ml���`Q�昷�;��O�S̯��O��R�>�}�Jwɑ��mq^���Z��o
~p�EI�DŢ7��M�������SI��C�2�YWT�N�I���#��
O�1 H4��\ԶP��@�^bG�A6~/h�N�K��'����"��Uo3�0��i�ZI9V~�9�(�<�Yk!fӁ�4B��e���%�jכ'>�4��?Hĉؓ��8�tˣw|�AbH*:�I��-FѴ�����M��.�����`�(S>��H���ϳ�� 3�m�j�=�r��.��fm9�B���!�+�nc�x��#�*����k�S�B�������ug�.U��?_�}$J���wB�`\��PL%���17���/���[�YS>n� 0^C2 hs��Vw���/l|���!��}#Vs�s�㐻W25��G���c��޷Y���LU��P�&�:����-|ԩX�z�Z��WM;W���*l��@;���Mc���x-s�������k�*��}��Y`}��� Mx3B�CU��_�:������N�%��WO^��b�*�z�oə�h�B�cNE��<���½׷N_�}�������ڑ�)^���L27oL��Bj�q��Ǒ�9��=(�}���s���=��D��	.<G����ׅ�!�8��t�v;ń2��Dc{C�-Q�g&#SN���Ō��_ -M
�㘑8]U����N�˳6���/E�`�G��f�eG�q���0C���g��2��JY�!>r�D�]
���~Ӷ�$x�H��C$c�pG%�]��� ��,��q���=5�f)a���1h*k^��G� >�s�bQ�E^��J����1�uYL�:�
���'��s�!�9q?j6\(�x}��c��"_�[C?i<=���)�v�e�Uhy�Q~�g��
]������F+9F�8�FƐ,�D��觬�B�.�1	�?O�y(�D��y�Y��"�P\��<�[s����c�U��ߙ�*Z?�H3R�C*Q�����-ȁ���*7�HN���^gA�또�s�����`U�D�mɩ�V�-����i
z�8G0�U�d��;�H���X�95��YE�*�y�Ħd�{|ej2}�� ��Nd��tw�"t�h7���"(�2�c�G��ɩMb�jj�t#a�G�����A&��!�Ԧ'�b�l(��E��4&2;��l�(>T靳�.N �+�F�����U�;��}�mv^�2�vd�Ϋ�%���N~���d��\��U���=�����3��]b^~?++�����3�1���8���
�i����d�H�K��Ѝgb���I �5���ҷ}+.�
&��!�25���Ք&Fa�7�0@�_����}�"Nl+�q���/��&qY���G�5�?(*�5fvD)TP�J�S�Ȉ��PW<R#>Y���W�l����<+V �BE����֜w��]�/؛.��ׂ��{�K�ޤ� EO8[+��Ӽ� �)+��4ro���T��`!��'��%�յ�::� cc�ٙ�M8��g��J�t-���k�ja]�~9:�k�W����t�+��$�]C�3��i�޹��F��=E5�Smi�?�ib�3����<ȯw|�����^�|�^D�7��[�]]j޻K	$Á�P��&(�MT��"�6r%O	�|ԯǳ'
�7-���;_���κ�9ME)zJ��������Zc�T�������7P�Lʀ�DyP	\�Hw2ny��S���J@��E(r�e��Wɾ�����s�R����E��36:duǩ�bĖ�*��~���i���}��;`''œ�§��Ξ���{�5���ɶ�%�Aj��K6��rባ����t��A�x��9��{�i�tCk���D�ٍ���a]��Q��_L3��|�wϥ��[Pp@�G�2
>�ʁE��F>�N�\Tzq�Ҋ� ���#`Ax��<)h��N`\���A�6���ċA���.	��-UȈ������ἐG=-�|xȤ��9�����-�q��[�?�~�!�v�;���;M����O-���Ѐ��3�HM=q�/{!c�� `���|�ү�*OK��0M�t���"*����_,�U/�������/�NM@�n��_g5�7Pi-,3�$�J��z�#r���H�#�'&l�ΰ��D�8U����2i,����V��{#8pB%���eq}�쉻�� k:PJ�Q�C\��𙦟�
���F�=cI��lv&�^��Ɍ��~�Նc���D��m����fWr�P�*�Ƅ�&�L�+��'U��¼�sB_�:`�ɯ	���S>���/Y��cG�vK�O� 8���>|Q~	�頳����p�� �.�k:	z	g �Wq��5r��k���?(�k���R����z�����=�bR3u�%H'v��~����]��'cd��;��֭��G,(y�����U������AVc�m��}�Y!�\�uL��P�b�;�Lyr��Q�"�T:u?��$`���^	�]T���WF�����1�[�����1����l<}<$�i�@2u����`��5��ù�p�\RII #��Xe��i\N���j�X�k?k�R���]���^�pa�x63 ��IYd��HI��&��!vy�o��֩����,�]1���K�}�������8����J���7����j�������u���+��u�$v	���F�eo����J��G+�9\��c��_*q��>����w
��S]f���٪|���(h8Q�D^�:������E�'�e �?�7�e	Pn���I*6�|s�W%�B4s����E<���Ĩp�S�w)��:��@5��솢���YPH2U$�&hh��;���k!tv|c���+�s�h�u��"�]+g��w�TQp��̔�=��k6�>ǡ�k,!�+TEWY �%�b�[/̀�������2&ȍX�*uY� �z-��K�h)6/Q��1���)��Kbldӡ6˟�@ַ��� /�IHۺP�gO��,���|���M�LQ;��7��� ��ޙ�-�x���o����V(Y���ܿ���S�)���i�D��}lY��*6���괷�Ľr���x����.��2S�]k<����G!�u:������AD�8S:"�Y��||�'��O���,$�Z�6C	��X�HD��)}!Hvʉ�5�@C�p��p{b�ň�H|�
��B�}AlJS»k/���^���_��#��}G]�&�6uN+�o~^��0��mQ���G%��[�ö�����r�~��C5�������ͪu��ֻ��%Ց�:�����J��UD}�06��=�[���EjɊ7O�]�F���?��u�-ř��k�V����s���I�<x)q�`"��{J����a.|%=:Ol34��+T
��zK��sN��<���2��g3��6�a��м��� �T�/��s���:}o�G�AE�cQ����o��i��i�`#���\�&W�=�h�/.��قIR@�Z���<�m�ݢ }����15�\�h&fk]�A�ۧ~'�ڑ�CKn[����H�x���� �Q�|�����S$�%�M���bgu~/�@*�3�&�rQZ���HL}�G.,>�g���栊LB�'%e�ԡ`+���X{�(�N�9"��U�~�3�W��?v���"wYz�dρ��w�BJ�̅_�&�7����k��pxMnй�9te^+����@��e��ȕ�o��M��\x|�iW�A�S�'���N-�B#Iq�+K���oY��WeL��OMD��\�<?�nu�>�)��y,�Τa�>w�t
:q��� ���6����!)���c���Q+�u%��p�-��̀��{��#]�p�iI���Ϋ�cR��b�6��ѩ��!��b���O+�b^��|ޭ�PP����*�B|�b��H�{>��}�S��.�Ć�^>O���m��`G1a��HĬy[�LAL�:��V��u% me��P��Tw)%AF�(,��`M 1��^�>�D���-ə��,]���ȩP�Y7���u���C�6�9��4B���>IƐE�v�;'H��2�.��+����j^���;cZ]�Łb�c�;�"��UT��G9������ij.T5�����'����j��k�98bu��o�"���ۮ��RLb@����Qv���,�$pCJ};x7�	6SN%�=�jw����$Z�h�t+��S�̇B/u�B�R�9��2��W9�t�t�.�TJx����)�6^�Q�;Z�i�%��͗e�m��1D��ߧ���ı���y	����#��px[I �� y������)$��4��8��-q�5�=fHz�z@�� �z;����#�ȫ�����jNF��K�I��7�)S�K�V��#���?�?�[����R>����g��9# g�'�~��_jZ;�V@1h�I7�?X��֧��H�Sr کh���*��"�Gb��\T
B���Pq����gek_��x�9�q���H<�iV^�~�_)�B�E�ANW�A�ːKU(N��Z�ﳂ�L
,�[5���P�Sr��N�Twʇ�[sq��D�λ��Ռ�0�����y^���Þ���4���T��U�h���w����>�{�[�c��W!@j�476�B��m�  �t�w�:�G�@B�&��TVXk�ͥr/��F�jВ�*�꩝>o�^�=PiN�cP�U^$�H��M����y������'8��ى��\k�W)�rw�~��+�(��K(ݸ�[��Ҫ��rYĄ�ԡ�&p��E���?άٝ�55��`�4=���O�hÞ���ϛ����лe?�K����/���M��,h�qB�w��5�oT��e�mq���8���k�j�`����BVU�3��e��e���C4�N8��&��p��+�Nd�Y���1��F�]�b��Q8g`}��lAx=,�AHng;Y>����G�Ga�5a��9jh֞�"���ڌ�bl�Es����rЮ�v�i��ٓ6�f��k�Qk�O҈���J'=�)8��Ԗ�.&n��y��&P�E����mc��]Z���x �~sc4���K�+0�LA�iz��Y��`|<���S^K��48�% �%���k,R�7&s�vx����)X
X��8��0D
�B�§���͈,ݒ��\P�T���R��I�`�U���i[`H"@=����S����}�q�=7�胵Fө�_�bo0kF�2���}u�ΘɁ~�G�B��6+��o�́sA�	.H� �|����"�k���;CRu�'�\��7G���
��#����Z�g~[��J�gyq6h��;�æ>�T}c��#�b��ێ�t��jɜ勷R�}���w��o��%s�`#�_�*J�u�>��us�P<[��#��X݄�Ћ��?��ce�G>vX&|A�1��-�!R��6,Pء��a8U�yY���ܡ�0ֈ�B3Ay��F�F�.ۣ�!����U�`��� 0`�W�Z� R�%ġ���孥8R�r���ͣ���E�����e�[4���؄~۰����/��]��f6�Nh��a���B<S�ݺ��z���w)�ЦgOսQ�!�hkN�ܨ����1�.���h�5���U�w4I-��7w}�(���sz����L�=!���r�Jf�å"xTe+^U�)�c��VcY��\O! �G�G�ZpDYY	��G�>�إD럜]�/���4�Z�\����UQa�i��_�F�B�Ǿ���$~FzXgв:����?�hU�J��#�`��YSk[�Ys���!�o�ꇻ��Џ{@T.)IU �|���g�~/��ij�Z@�iK� ��҅M��X�"M ��$&�o�O�1�8�*�܎��9% 1Fi��5Ź����qҹѻ �I���'��u<لc�- . �K��1I~Ħ.�A��?{�0�e�/��������qv�� H�4���v���Q��YHO�����`!Pe��'��st��^�^����GQ�����L�9Ro.��~�^�T@Ot���qrDـ�[6F&��j_ܜc�����P=l3�.���a���A�]E+�dN��޼�w�*�y��`�t�I"Y�v�W��Hhv��%�Ĳ�������-"�/ߡ{�A�b�%>Lfd�C|^f��]F��V�OB�/�U��,�:{L��k˂���W:@�7:���PÖ9�}�h<��@�6,u���F;M���[鈈d��H���m��Yq3��Ж jȣ�����+����ێ+�p�&�_�M[�(o����@G�=-�d�U�����*�pu����h��XV֦�4E���)���8ڮ���[.I�kdP��J��<�~b���k %x��{���v݅��\�~�(�\���;+�j�ix�;_�8o&���FK��� .3کB<�W�-һ�t� 6o�p1�i��޷�g��>�Fw�<\�>z�Z+G���s�|�|�e��Q�z�����{F�=����0m�B05�<�$���k��t�8����m[�%uY
l�$����J���� �u]B$i4Ch�E�1��]�_эCf�lcs�6�#\��%Ej�b���cQ��he(,�=��	�����1O37Ḻ��Yy|��wмE����V䤑�t��N0�a�J3?�������q8蓻֫��v\;��mE��0�H��?��-X{��
�����b�]@OB�����~���d�QLu�>X�f�����P���J~F��B-6��[��#]߳�1�oRl+|Y�o$�O�4��?
��J��������9�B�$���ʯ��V���F�Cɬh�4Pf�ϵ� ��D8�<�܄E{�;�k�]��e��d�A%`�=No�#ɉ��/6@#_��O]���4���(���F��Z0�Q��[ZwIss�d�O �)Ӿw��}bn1"�{vxwU��ŷ� (A_�i�#�m�������ӣ�ϲ'b���v�Iv�^N�ޘci@rM,�#n&s���6&w{'8a��{�Z*�/tAH%-q�,�h����϶�x���󚹯ߍ����#��=J��}Ύg³%F�zo'rC����U�d|$��V^�N����_��ZJ=��=�KlZ1�]r��?vtXc��OqYh1�e�:n��8�I���\Hi�.�{�9���[�NS<���w��o�ꮎ��Vۼ[3����R�?��\!�[8-bw�D����C���_���;huǼq������ro�C;F5��Ng���V�.|�"�D(\�ߧ�u���� H��y��1r<��Rֆ�]�֞��k�T�s�X�YRgU_ʡje�QX-� �4-#��u0J��+ɮC/(>�G�6a-4h˳F��o猙sՐ��ǒ9u�X'+&]�!��K%��~��},�m��"*�����c�·f*1u�ۭ�oo��}���yT��0"%�T�~�]��
��VTdÞ�(!@��k���1{�<��,��rY�5�=�
�V���l�U��"��E:����H���z绡1�w�N4ܵ��"�f��?���=�7�{6��*��D����VZI<U���i�s�W�3�c�ck���*�6]>�7!E?b�3ސ�d�lV���&x'�Y"�fQo��;W��۝�[<�em�y�&��/ʸ��'q��%���I���6���;������r�d����I3���^K��i^&�ԇ�o(�D�{Q~@e��W�*�	���)���D|����o��uQ�D.
��"��\ԁ��큮��[�1IA
���v�� :���<F�$�I�h���S�(��Y�M��Մ<��F,��\�g��ݒo��T.����w߄�LZ^U��5��c�w�
�DN�E��������A;Đ���>�����s��t��c�]q�>p�!aV�U`a0�b�v,�m:v�ٻ����軱W�������n���|�Z^�^���_�t�/���E��`��N��׎��؞_r��j���v�2?bŠ�D�u�� ѐDV�*a���!m�i���L�H��!�a3��/���ߓ�k�;(`W+ k���K��ETѿyv�����P��`���}+暘7<Ѩye�cS����P��*�$E���Cμ������\��ߙX��K+�*�0ȅ0C�s�V���'����J)f������4�՝~& J�جcILZ����6ɲ��H�Z�qD��4[�,�����Q:�iN�z�A�n�=�3e��4����m���?b=8�P�w���=Zl�E��$�ܮ��=��y=.5�/���6��b�J��#?ʀjN��ϳ�?���ęт3����ƨ��c�Ҳ��dL���HĜ��l�9Gۙs+*�8��a8Z��\8}�)�o�&`�r�R�	?n2�dWR�{�|Ya�Gr)|�Y>u��^��+YK�b,-���i�gRj<�{����]8���#�~�=� -��V�T�����8=3̴�.;��U:�;;�n�ii7%���Cд6�xʶ���m]���%T�]�����������b��":O�JV~/�^����=qЂн��	�Ш��olii;%�o�VVb��O���}n����=�Hcy��24ifap��B<���y��m��5/���v�5E�Egݾ�~��Ǔ���Ӣf�����{�&�Iz��N!T���0�|�${�Ϧ�w�`tŹ�pB�����4n�5��W�
C.2��r �s��Ɇ`0�JW�:rajo��E"���ÃR��B���=G���'Ku�ʋP�!s쳚8�J�P��>����Z{4�?6�[�{8V�����P�FVRTt�������y���5�ʲ�^1&HĞ���E}�-I�;,��A�S�%�P��U��v������M����d�D����%�	��k_�:{��TAoz�;�j�2 �����NB�w�O��lx2�Gd��1���b�A���H���]<Rw�>��#%|�����&O��D��|!f�ц���&gٸ扄f~�_�K�j������6Zy���:����̝Ij3�M�ojz|��b��6�P
�5c���a�}:�ڣ&��=qdiS��Ew'?�߅�>|�g"ͺ��n�Đ����U�� �ꚴk	�y���.]�^ň�������k��5t���(�ѝ2��4G�]�8xBa��2�7����<_Z|���ҍ1�;��u�n���}k��rU?�\�r�����ҍ�8<�/���7�7Z�M�G�$_3E�����N� A������hu���u�Z�K��̥fb�F�Qe��lk7�Y�7�[+!��u8����,�Wi�
i�h���Y~B�ţZ�F���N��@�}�/�o�րN-��aG��)��.ua���mRwҿ_��ϊSURrV�^�G�o�AB��~.���,J��vtk�ɛ�Ƿ�ht�ݦ�����ꕃ�c��6�H�M���\L ~�C�b����_C'C}ɤ:�W��TۺW�8�����A=k���#\��d�O�+9P��}�����?�{��D  I�iO0-�n/aX��׶~]>u�keo�H��B} ��ͳ4�Z��l��)@�5��.���I�M����
^,�q(��Bc���?�);�cOkQ1��x7��8W	5��/�&҅l�9|��:��?j�Ǧ[TpW"x��/}v��w)�����9��������썿Ͱ��qp�h���)!�="/ap�.5��GL��(�V�ty�O�{&�)J!ֆ��7=Y�V̧���MH���:��|A��0�+�vq�pM{O����Q�w��t	�]kr,��6�C��3c�ɑ˷�l=9e�㟔�}u�A��R�ѦZ�ˈ�[�_�#Օ��u��xw(�\,=::��m�h���)!qk<"�ی�/��.;�O�2ȏ���Y_�~U��~�}�ҹ j>�K��&�v���X�1�����w������g��J���������67�-�k��$)!y!c�?��7����9
�����]�����C�	j�����{
R/��]}�
�Y���K�^Y�y�5!��R)��A�*�����P�CH���g�T�,�&c��{t0L/D�r�(����<$Ѱ\���.��i���Ɋ��&!�8\��+�J��]9�˔�M "�=�a+����ԗ�u�h�I������8J~�����i3V���ÀM�F��S��FuA�L�x06Q����p	r�J�-�����Q0�%ay]��U`�?~arxPV��'V>َ��,p2FI$�y��dt]�T҂�	���7��� �!��P?Y�~Hs�	�.�{�ﰊ�wy��?#��3��Kc��|s#��#�����N~{.9���
.�H5X�|�f������ ���j0�#"�O������ó��vo_�q��p!�EB���ߓ�**j^�Pi+�Rffx1��%���I����n^#��}˝��O��"���!HܧI��r"��_����W���Q!�PRS�SW�Exxۯ�6�P���|�2��*�V�8ސ��-?�|_̶��o���OC�b�H�Љ�O��ϓ�5K��e#�#��;��!�7Ϫ��h�����zK��k.�&��*��U̾0�d��gƓ�[���%�j�7q��R�����Ó3����L� R?/Vh��kf���jL�Ui��L"�n��~�v!�j���0�.��e�����q��A�U�4@a���{R�E��D�۩���M!'�$�1�9N=����YVZej>��±��3�("�����+�����p~ޱ�r�`a�D6wV�e�D�IN6b�%��+*�������!+�9���n��
��$4pOfkr�n�m�Ld�zQ��$��q.b&�o�Mv���Ѩ��,�^�������q
�r�I��a���i������y�cG�ŏLt��˧���R��*�!b�G���	$�کO�^�u�1��Q��8Zݫ*F�z�Gp5��C����*��W_d�hӪ�F��8<�Ir�p[wf�:o`9�RI��$V��g����<){��i"~(ґ������Z_�����-�l��SH���7��Q&c륲Ȣ�Ai;q���W���{��oqp�T�]	��Ym)%�o�ӿ[�ZO��TB8�9o
C�\��zk^�7����y�@����٥R���/�F��u/��#��NA�N
eٲI�/Y�����d�
��B3�
��'�}7��p�~"Ih�1%.3`+���D� ��]٫���BXF�;�,;�,�����R�/�;��".�6"��ڊ���b�L���?�^66c��|��$o8�ҳ����^8"83�����,����i�o�q؇ڔ��}�|Φ���.�z:�ɽ_A�S��B�+T:�3��E�����8�M�[h�AJ A0�����}5�664��΂���xMZ+�X~���sQP�g�u[�X�=T��aE��_μ@v�I�g��Xi�F��� �#V�����^���ҷRDF7{�z���AF��˕�2-z��au\z��ӽ�6�����=�<�.�}d�fk��)�*�-��;�N��1�9�g��m3:����wHz�mE������!����O��yYu�B��˰�HV�ab'��J���6�T�5<?�Xv�_�(ZY�.x��<N�k��G&IPV?A��2eZ?�*�L��h��5
�V������"��͞3��p�� c.k�{x�l�H[�~���|�GPLY�P/
�H�/����b�!|!��Ps,'UF_I|G��q,�r�Q�.ʕG�UU�7�����`��u��^$U���BP�������K��9��p��1�:a� �j�=�@*e�;�R��˓��5i(���l]e��9B�cqC�$[�vy#7�U:��V�mM�n�D�"�h����#���ez�����	���7{����J�«����N��cG3Z��=���8�ș�����c���Vt��D���3�?�c�qج��-���MS�t�T��~Z��I&����$2L8K��p�7*6:3��:9~�k�X��3�꽹�$\�2�X�����ߐ=������57]��W�S���U��������6C�Aq|?�5�`t{��hF��=���v�dL�!���(��.�gg���J> �[A0ؔs�^�	j�vژ�pBz�[P�_/9-\l�ܲ�X���y�E0��0��.Ż�����~��y�����.�1������,p��8\�w��4Q$�f�U۹{��|��O�)�$�<L�&��q��̔�ԊM��'�!Cd� �w��H/��� -��b�H#�Hd5t$�zi�����Pχg~��w��=����y�vT�<{�35�eR�e~
m�;�Yp3��;m((���;9��~I�ϵiEyWW�%1Y�GU��1����@y+�H�@��CJ	�ȝ�F��3l_ө���EZ!��?����/��9��-�#��l%T�!fJ?v~^D��3��.���+:t�	魩�(�}���zU��p!)-ͯ��2	��] oALЍ��o�S3V�%'"�]�D���H��Y�>5iϝ���F��
�H𡸭�H�^�s�h���1��Z��_4�mN2���7x���@�E��E嬨�Z��� ��0stj���I�1�͖��?$c�|��j�l�	�;�I;%�P#z��gs>�n�D@�<A�h��G�C��q�ᇥ���ux���)*hԈ��춇G@�Nl�b�cԻ��_�a!t"Z)��������O��'rץXW��#]�{ߌ8 @ߠՄ�-�mr�Z<��X�YP��\�U��bBZ#-bFf)\���AQEųmGq�ⶒ*��H��Z;r����� �٣��:���r�b������6(�>��A>1�4Pb�`o�y��\kV�V�G�T�w#���Q��B#P�x.��q�Z�c���-Ex!�l�F��\w���⬩�8h�і�(u�J?���P��OO�F�c�)���r�̩���Ó�Lߥ�G?×L��S|�:��Յ��&�!o��hZ�V�r)����P��H�̙Or���{�
�
��8eq�U��b�?w�����y�vj�%�g���^���}O���]KKD�,�sW�� �ׂ/���z����kok�x��I���SD��iA�<	qmY���֋!��\Q��225t������O��m��"%���)���.rv����Ƅ-��#��ڹt�@9�~X����y�N{��O�Q˒*� ���[hd�Ŋ�|��~V]w~�A�}sϳ�!��ׂKP ��yfb%��\Î�ŝ렆V@[-,j�R����uŧ���C������4��YX [&�����	�=��z�@5l�c1���z�FC�n(�����i����[q>4�ޥ���ċ򿭷��uƺ�tїg�Qt.��\L#��%��U��'�}�G�����;�x��/��ݚ7����M����I�%��jG�&��5�֋���wBQp %"-�at���*���ɳ봭9��8R����y8��CcE'��85�]�����#��=��Wl�ŔY�^���I����`6?�o�lg1�����EEF��z��m�6�C�%�������_��RV�����*-�oo���>�l/z{�5�x�P�7�����o�ɴ~�������c6��＼�F������V�hi��-uh�&��Q�ه;����k���$6mK?�3�-T����� F�PJg���(Ǭ�ލ��yҘ����U?!e~"�cY�Tmv��g��06�����t;�&RN�6C�s�6�Kfj�I�Rs���#ىuh��6��P1
����K]{m��S���,��C�V�rNq#�<�Z����o�n����+����J�^���G����j����,���DObiC� �6�TU!~<2���zd�¥H~<��m�ڀv	�����^���Q,�dc{���|2cy'�������ש�~퐻<9����eqQ�67�i�=,�`5��И\T��V��������L���n�h������W���x9WսY�2���c�<�ϘlB���+�p?ft��6�#�D�����Ű���ҌZ$j�o�@,���ؚ[f��*~��d�a�f�H>b˨'�M}�.r����P7&0bl��l3�y�]����8B��4�1���p�6	�$�<����	���r�rs����~s�вhv�Fd>�������֧֭��}���Q�����6e�@t~`����L(����ؒ��5���bL�n�[{kQ���lf�n��ym�rp�֎f���\;99���(��l^ʞ���;�:��蟇�]J 𵻅^�AҚj��9T���8\�3�����'1Kj��J��	���&]�͂FQW����+�#ke���)��ogV&�B��th��c^!�����+��j� qww����N�����Awww���!����߿��p`�7����U�z�p�.�ۜ��x7%+B����T�K�������+)��(���^����n�b�w+n��=wmw��8}����bY^��!�YbI�o��3�������P� ��V{�Jj�v ל)pJa�nGQ��>��R�d<����,b(K�o����ܮ]	)��٥���.b�~w3��3]o���m��O��=f�WI+*�/���r>���$���"��N�d�"7�;vV�uŗ�z���a�V��=$��P�^B�?��Z�A��>P�Z7�+�Lϙ�8�;{����;�8�$�'`?���Q�_>�)��T�6k|���"S�kF���,<��Ltnĥ��4([C!}$�--�Vsxk��r�%�o;��ۃ��3Վ�i�n�1��&��'P�1�F��L��yfc���-N",.m^%v!�p�$f��F�}���kO7�(�+��YA�������k���S�e������]�Hiii������W..�PT0� ⮩�f�M8��� ���d���8x���)� %ā]�_�~�ӖQ�yv�[�BV��V���	M�-���o�x�D����lxPlu�����@JS��n�DPz�++H_���̙�M|}˫k2�}�D%����)�#�7I"�s'�;NF��)!�'K�IX=�/IB��م�Ӛ���QĂź���T���>p����.��K��( ��=���pmm-���Wc��C'D`l���G[�JT����Lh��7��/?�.|,�W�pF��`_ �D�>o�����0�4��M���#��7��zj�{�޵4%�)tdki�]�>�
���Er�d��:Ҥ�y��[Q[7T=�I��<^H�c���YC��8#�����,������"'�<Pj�B|V�~�Z��؛ӑM����F��x�8b;����P6��ï4v��H�V�y��Pa�---����u	!O��P����5-���I6X����-��yvV��e�!�QN9\�@��i�*Y�!|�QJ-����_���[�X�@T�T�`g�,^F�
,z���%FL�{}�=�W:��{s�l�d�r�a�n��تL<Ƽh�������#��b�����0H?��n]0y��eMt�i����7ڧљ���Ȥ�L~�3D��',�ۡ��n�k
��P���?<�W�6��iI����[Z���pp`�HΤ"�*+������P:[_)�& ����rx��%��￪����o�k��o�uF��PLMM�ă��h��tf+.��!���c�=N_^�ir&�����EH%��B>h�5��I0t�sA�=�u��DB�cB�qm.�/h�oũ�7��K���SsR}�^ę�U�c�Ѳ��А�u����uБ�����7u�V�������0Q bZ or- ����I2r9u5ҥ��sf���ë�����c	
���Y=�/^?4���F��]������F?5���j�U�����'��������tE��1!�K��J=t����M�eԯt��< �ZU�V�:��^$B�sև��L�[��@G�|E�|���/i��}�Η��_���*��JuA8x�T����(nN�/��y�S3\jX$Z ����e��i HD�V��Aa#��K�R���즥T���j�I��cj��sd�y?�&F���IJX_�'v�wU�W<�[rj�,KPLFl�i�a[{��j`H� �0�D+�X��n<�ʽ���"�d��k�O]y9��:���9�ȱ��n�v���T�r��_�x��_�����
�p��t�ܬ�d��<P�OQ�P5ăA5^yՈ�:�!ۇ���j��;p����{T���t���B߱�A��)�s�lo��r��Te�F ���b,h����r��Jħ����zT����:�� t��X��i#���&38�:ː�	�n�Eɐ=lp"�L�� �"��)4��=�����
c� ���A�6��[�1��m�����z�ֽ�{����.w�L���I��k���I5� M��T�������K|>I���d�	o�J���圁�c%C�Kio����y���N�����zF�W��Ӽ �!ˊ���8��<k0���<`����Q��ǖ5鉫R�D]����_!�s��[�8Ȝ/;������	<e���2��N�Jt�:a��V�&��+4��D������S�p�L!�έ�Ǽ�Z�G�Q�q�b^�0<.��2F������8na.�ta}nN9�,rwB���2�)J��5�g��Ks��كU/
Es;�q�k�4",�����%/9��ӗ�&�d�8�b��t��V��ݥ(_���{�K�B������j�,mP3�@��b��- 7KeFFщ��
Z�v�Ŝ��ضJ������!.�3�ʿ�iyԢb`g5� ������J��_�o�$E��L�׼"�[z�OUj�n����߫Ϙ�t"��I����%��;�Y�@u��KG�SOG�1ăVfNKF�SF��Կ�pȍ��Bf��Ahtn%Q��9���D
��R�:��X�]n������`$zm���|g����ؾ�q�K�̄��({��@�iY0F�$
��=�Zi3�qE�,L7���|7z���zј�f���c�znIL��3\F*�Z���9!#Z<n:n��9�9&〪9s��/I0�g.x�NȤx����*0e�b ޺�ĖT8�L��\A�ʈ�(�g0�������FA�Q�a	ѫ	�F���y�e����k<���ۨs����@]��㳻hA��$û��fdk���~���,����+S�R�4�:���M��ú"z02�q<�k�v�ʑ�H���U����p����iLI��Vj7�;���cI�bs7|5�?��*j�\j�ײ�T:�j��\͌L4̇�Q�N\������/��k�`;1�����4 �G�B�g"f����.@AVhͥs���r�=���G�?ت2����S�x"$���h<$��Os|��nQ�{ �x��Kg5�b��D�ڬД��xJׇ�1"M�C�ʬ_��]c�T���`�V\ōy����*B���9+�dqW��KR<�i������r]x4Uw��k��}�FNb��%�qt:6|*��P�{�O�s|�LP,�� FƉQ�La�y�&U-��u���@���Ȅ���p�n^]G��&{VZ02J�%�)(0Qc�:fb�ķ���@�i7V���3�u��q1��\zؾn�Q{\�T��b�Ϣ?P��8�܈#�D����˿�W�����u�tu�S�B�i%D�l����P~�Kt	�iRF� D�1�-):0|� dpa�a��w�U]W,l!�<���
��F�H2��U.��,�r7u���.I�c���,�pV�"G�ee0)0��GA��Da�|����Ad�%����r�dɄ3��p#�#㇀&��
o��1��[^���U
�f���c0�)�L�A�ą�de�(�ŉ5�~�CG�Gxf�Z�#��r�D���ķ�F�S�N��jG>f$S�WF�TP����a�_W4I�*�׻j:�yA������`�j� t�$F�1�Z��ʣ��x�����8M���g�M)e�e�sHR�Jit��cR�� h@����Kz�u%��+���� !�����b >��H��(�`-\D�b0*�(yT��1&������a�����.c��7���v,_4�"�����߽�ĉ0)'d�h��_������H����R���~��=�+��H��T�	��4�~DZ���3�F�����뿘��z��H����{%0�1Za�p�t_OЇr�>g"�[�6�K.�*���+�FNl����q���k(5��F.�豮%�0'��f��Β���&�C����G��p9g�`5̨�gnFR�	��(���;U&}>G����1h�	����tp�b��!2��3�v�x���G��ߡN?�P�-|�ߙhK@;� ��33��<6V<Q�#�_Q	�8QX2�e��%ѝ/V� X>�:�+����o�6h�Nk�=F�YnFt�AKC�i�J����ލ&��Z����rRG�x0��*Ng�ܛk����� <M��P~M@��+�\q0j]�jG\A��=HDv9l����-�m��i;ziZ&GT)�;n.*g۝�ߓ4�ɐ�(���D���	��D��|�E�o�"���C�՜"��)��NF��|�q�|3Q{�(��=�q,X��\�f�s#S���}�MW�	]�:�zO��ޜ�Z�����A4$j�%u��wPh���U�������J?�'�*XPvH�Z�H�̱Mw���L�V�� �&��F��K�*Z�x�j*T�o_ݥ?������cO��
?(т�^6ph���5B�W8"~ȬI�'P�<o��ʱ~3M��)���؃ �1۠|5M #�n�r1��k0B�W(�x]�χJ�Z�͟��p�v0t������� �}��H�Zi�����=H��=>�( �tQ�lCX�W^�����L�d�gb]R%��i���}��O�d��Wa
;����Z&���1/^)��kBD$�N����Iq��gߐ�ˢ:�{�=M����&���%%�����4���9޶M�(8YZ�Zb;�|1�9hfv�G,}���4�<i�ѐ����m~]��M�g�oĕ!^}^e�%Q��$��z�!Ѽ�&G��,��H���F�
K��ϻ�)s��HO_H�3~��c��bj��̛`�]��	Vz|
B�����t%b��詫Q�������ҏZ�b����g6ܒ@�i�=�I<$u��X	��v�R�6��Y��
S����%�O�Jԋ�
��g�/��|��]�/�g\m�I�Rc؟�YJԋ�@��!�؍;�E~���i��L!ar����,��x�o�7�E8r���<6">]��_�BS��&�	6�w����Q��]e�E���Ѩ�E��������� �H��������m1<����ƺ[���Ӥe�g��	�� Z�d���$2
�J���Ot ��NCTj%��,g {P�ɤ�Xs���Y��A��\����Ru �`����˕��/cGI�tE�f�TE��A8:��*Q6�y+�|����P�j�q@�\n7���P�J.v"�k����v�R�p�D�Q&���hMoQ.��fQ9�X�M)rتt$S"�n2��$��եwmSm�Q-)�^G㾌nl��4X l6�ئ�l]=�����rbS*�S���)�#���8���-�x�qkS��~vFj��t��(�fl�v�6�y,�b:���f00�X�,�k�XLţş@<6 KE�&��6E��hOe��z݅�	��̟���<MF���T�V�y��)�%�5$�����u��Q�k�D�	o&�����.=�p ��@��PIϞ
E�i�P�U?�&��2��S�U ��!����<�� O�q �Te�wlᖽ�ܙ�״���>0�u��g=��ns��BP��D�OB��|����<��*�@'��݉f"�A��t���+\�6��뤦LCm]M!ߐ(�35���2,�MT�������VL��?3������S�YI �G�_>�f�76� j�K�� �3�DW�L+a���C�q��,=$����_߻Q�Veqb"��k������n@o<��7e�$f���~�'��I�tN�	$��D���޾没��}r`��&�1tR($q����-*�����0(�G㏃�d�Q?$\���7X5Y���؇��fm!L�8	~�\��9V��Da~f�� L����ig�s����=���x� �84x8R��.�*�O'�OP��_M��HK���^u��x���x���L��X��1ߥϚ��$ܻ��wާ�ʧU�[]�T̎��j�G�u�z
�E��3v���9igeW����5����z=��������n$�X��N��8d�kqOqH�����m%�|,{F�������'�c���[�)n�]�Wm�Z·� FN!-_���X2�|pdCu�ob^��}�RfDy�>j� �JX5�\����*Q�Z��?��"�|��^ �:w�~�~�z�s�|D'Gf<剜i�����z�6�y[����6�"tw��p*�D8����y;E{��~'��ZC��̮Y׍�=C��U��ˢe'닮��ʯ����"��A���$� ��{~D��	Xr�8�L�\`�S�̎�c�؊�Gg��<̊����P� flL�jʹ���*��Oµa��+OȈ��T>=�±S���Ny�:��[��X����~�yC7><��{�h���:�2��26웈�Yk�x�W���l��j���N#v���=bܾ_1��wR���۟�S\k���||L��o��I���v�/���j�{ ����z>�,���D ���e'�v�G\8`k+�(�P��'��h0�W�+̤�j�*�qêSu�h�cu13*�D:�N'Z��!���A��E`���O�5C%���Ꟙ�{�z���Y&���P����?���wF=�o[n��7Y�p5ԓ�U���`��b�_F�U[�`��3ǩ<M��f8��](��c2r@t �0����.N��X_��_�Î�*����Nn��ȇX�ݜ��Y�������&�P�S��u;���s�I�k ,8ks)j���������}� i�~#o�g��~�4��]{=�*�Ki� �!8����=�1b��}�1Sg�2U+P2��L�˿C�5��`vu��� Zv8"T[�r%qW˝�D5L���D'�4�~6�,<T%�\D^^�h��o�1��#)w&�*jl#}%�����rp�XA������O^>�����y��ŤL�e�B���#}����2�=�}<��eḦp����A�Їf?\թC��0���4��3�-zN�o�Xy���rw��e��D�нM�#w����{m���_%�I��%���j5�}��)�9���6abT���vD'�i%A��0��k%}�wT��Ɗ͉���W� ���)dF������4�t��� W�0�=�Jj�\�,-G�Կ�Z	~�2�Q���P�P�iX$̧5�E$�8�b�R��1�7eh\r�+�!g���}�8�429x\˦�x[~�E��I�ؾ�g��8��`�������ha^7bFvqI��;:�0���N�lޱ^�o��?Еh(R��L��ȫ35C�t{�����I��+I�0zu9qII�²�-�e��fh1��H��`֩�d,�����_m��((ŵ�|p��ߙǧ��� ����Vx���[�����	[��b�������+W��ܨba)��A[�^�۸8�Z�"�������Xm��*B}�3Rb���y��z!N�B����%�)ma$��Cp���8g�\��(����'Vk���R	��k��R�y|��#(�$j4�Z�_�N�9)}}�;�+�#;��y(�Z�7`�%~�m�4y�Q�ɳ:K��\(��ݳ��!�H�6�}�ǚ��X`����.�G��1����׻ƒM��	��0!5?Tt$/7�eև2ɋ+jTd&&�y�ާ���5�gw�h{`�݅�\m�l@�T�:����Z�U�HIea���3;�M"����tеƏՌkQ��L�0*��1�6�"+q5H,�	f��ě��:7h��iE��η4;'���\���C`m<���T��%35gx�h�B<�d�P�i�lm�\�y�� KI��Et咿P�"A���l�2�t�����im9�J�`��6�߈y'_ڹS0@�-���7QRhԻP�\^د^�v�f"�>�a$u��-�	�[�[9G=���Z�=a��Ɏ���L�2���C�ZX�G�`�	���@�1���Y�K���S���������t�.���2�8FM��N��g�#�5^.��ِH���S0�*�ϯD��N�H2��ޯ&y����q��z�]%���򢍮�M<�Se����YJ
�;���
���V���g�k�1���_w9o#����߶"�>�/Mt��$�	q��F�|`�W<Y���s�34\��7���6��]���W�Xъ������HH�^�*5��C�ܭ�2���	iB~7m��N�Y�$��E��j��so�P"j܇�K�Z��ԩ���̣�`3gy�ܶK��� �� �ъ�6��g+0���o���t���'> 7�c��Su�����:��CƯ�������_�}V_���Hv�Db�䇪�lu9+�lXN>ZyE"Q�|�$6P��HBl� .���bwN�Xj�'	}���Fo>�]�:�/1qM�Bc�1=AX����l�~��
��N��wu��e�b�ԏ"e�}��n�,�5�� n��b���nwt*�(2���e��/ԅ�
�f��)�i�;�{�60�·��[+��?<6F?���o�~�ɫw2���޵�A�)KA���e��S��_R.#p��6���` �'?Iۦ}�.3�'�;!�"i��_��;�/fq����9E'ey�d�Fr��!�e�S_�D��@�����zW�ER�{>�).)u���u�B�*��w�������[?�����6;ﾛ	�o�����&s��>I��(�M��B��A��~M<D�↦�bq�W$�N�������<�j��M?��,�m����|\��G�OV'ey�[v&�p!$�r8��5�0g�����䣫�����L�P��cl��nv�;���}B��p'h5��C���ˊ@���R�j��O�|4���Z��xL��xx����^�t���.�`3Z��IȦ�.rsRI(
σQ���ri��;����1KfH5�uFEB2�̠w#:4xg����Y|��fJ'�j����&�h�����e�.T���D�.2�x���a�u�%q������fH���D�G��\�'�#�� ���+�+׻���_v-B�Eļ����k�[]v_���9���-��m�*Óf�׳�%��K��Z��ݰoy&�N S�n2g���<R�/4�]['��v:�q#`�?��L�*؎<	����V?hs�4%z{��t���}����eQ����)�;O�>�zbR[O+Ҫi��3=�9z�u?J��d-�AR�W+�,<ؖ����9Ӱ'���Q�Y��9�b��?Y���
��	�'��Đy��Y�v}�X��',b��o�x��p]��	�O��X�ҟQZ-y����<ʵycxU�T(@A�0h)�����0�@yh-[����%D3�V�r���3HP���S��ŷE��#��FtϾ�;!L*,��m&U�i;� +�B<� /��H?�l�`�Y�K����p��8�=���v�Z
�b��mt�&��O��Y���r���]?�1��o�w���l��ؐp����L��V`��d��%餓�&�������T?.$�z�F0C��e�by��p��$���F_�X%ϙ�����������	�?5���ml�z�������xU��~�������ȼ��u����g�����ޥ
�,f����jsU"o}�LGٓ}�^�X�P�x���hM�0�4B �cS1��o�s���ݐ��sd%��Yzl�ģ���9�*`�kj�kNU9<]	�u}��o��B=�+>z�Fr��_l0�v� ,�y]�?�Ѷ�wm��-!쌡Y��[����3��������B���t3�K7���#�� !-ºK!�#8�s�*���Jp�ۗ��dO�a[��[���" ������ǄşC�yQ
��<#������X�����I9-�ܘ+��Ȇ.Wz������D��H�N�7HZDW-QK0�.̊O>ϻ���Pt�Ȑ��B\6z�՘�D|po	�X�'J)Ϭ��1�svTӣV腀~��K���S�NB�83q�zJ�ז��گ�á��r�o�Q���hͧ�|&��0@��S�j���|�{�\'���Y� _9�B�O�P����+���[Ԟ��gš�u��BT}_� �J��A���O�X/��)�p
X��% ݂�	�� �B��
ε�8�s�gF�I"�S�j�w��j�q��?�E�(7kOO�1�m��`m-���K��<=�ѣ�t,��8��?n�zQ�Zʙq�ˌx��A��z���=�E�H� r�[�(t�7��V��K�M_��P��(��ة ��c���x����$L!�D�j/������#��'!킣]�]R0��^9H�*l���ӽ(�F%��'�:��֭�Rf�C�r���4@F�S�_>>��BtU��t�s�Dwe�ި%�������T�!	�d�3sm	���(z�?�G���R����z?X>��0E����6��7����C[�;0��u�����=����Pb2�����1e;> x���p՝��Ƚ1f�q%��p����'ȫ��b'�J��	�>F$/�Fm���P�ˑq�_����HQ�A�i��V.�]�-?�*�r���Q5�����a���c�K v��^��~DS#;�/��(��~�����Ϝ���&e������\��R���݋����^�z����jOvS�F�]h��-a*/��T�J�eFc
N���~/ˑ~�Z%�s1�L��/(R�í���н��Q\���ҝ�u�uT��ܷ P�;1�=|��5�U�L2b��{L��$������!.9���!+(���Z�R�� N�-��S�`�[���^N�;L,8S�\X��s��0�JG#(t��ޜ��ޗ0C��O��$<���\]5u!��i��=)%��L�͹�:��z�t6w(lW�b�Yn{52�L�f�4����
�.�8�ղ;��g �:f�d���r�m�o�V�ݜ�'�	����:���6_�\i
�����b]p�~
 ���;j��,.�������f�S��b�\u��:����Nl}��[��tE��jČ�{/�f8��)b��EA&���@ļT6�axXퟔ6� aRvgjtV�H&�+�K3o;!��Nkz�1����Tk����oN�P����7���uIl�,����̮�i8{z��K�'�U��y�/����,|E7z������zp"�?��z�U���k���|֞wBp�23y��� ɶF�2�(x�N�[�@B��LM�-�K����4!2�����e�h�W����G{پ2�ha\kĎ_T�Mힻ���d�X�7t$�́�__�c�rÚ��P����ƀ7��Yϓ��y�0|�> ��a -�s_��ȭ��b]݂S葩��|81B��C�5����֤:>�K��,GR;>�6/d'�E���(�|�T���^7���{:+����L}�i�.���ʟ̸VF����{�"��v	��_]�z�~K��Z�){ի+Q��'A||���l�/�2�D�9��'H�;��;���`4q������p.���$:V�ʫ.�� ԝ=�pei����i3�m�L���JHAǞ��K~�ֻ� �����,��T4OD�N"ʹ*V���5q��/z2�+�����TO��D����}F
6�I���/������l��p�D�4W�Xѳw�{V0t�|�E3 ��ٺ��]�D�<��g7�I�(V2|�z�[���m���M� FӼ�д\�]�}%5�N��ams����֓��?����r�E���k�#x^�<�5����
ѧ�4�"8��^u�l�����4]H�$.��Y�?�ŌUNT�r�IEq����Y���}�n k�<�����^�W	�w��ED"x��-��ʬ�����K���ZV1oj�0=;�{�����Qz�͚R�c%�ps��VX��5��L�W��L�i��������D�rP�R�3��&��]&|������b�HQML�0#Em�p�zԩ)���Д&m�Ek��B�)V$Sv|7��iҸ԰]i٨�aI���p�D�&0J;��>�P�ɂ?wo`�-��?��|���?O>��R�y���>#���L|�Q�D+���ei���.^$t{��&.S�֛b�;A��`��#YƷc���A\�8���7njp`O��ֻ���9�H�]�O-*ϯ�a�Ajj�#b��������@i�۰R�`�Ǫ�i��˭Xy��
��@D禉c�1C�ޘ�m�+��[� �ǫ���CTw�x?���i�AK�~*��02�3����T�Ԍf͡}��tz]&��ސ �h�n�}�J=8�;-mF& Rc���B�H@<�1�,uGS�O�c�E� �6��Ƌ�tN4��{�.Q``��z�iP�Tfjڮg��JKd�ع���u^.�t;�y2����4��e�A�u\/������3a3a@�I�b��V��Q�2�=�{���������f�>����`��[~s%�[�,�//0���V��~X�8X�v"|�a�*ணf��_��6�	Z�HZdqrO�?�n�-�I�w��6�/u��!�6�j��е�	�J{ �q=-�L�B��t�W��;n#��f�y�rÿ���ĿR�T��v�ۮm��O��=)�R�PN^�������f����z-��nC���B^��0���#����Ķ	e������שW�j�e�uX$�[�s�ß�S'��g� ����<��02e߇_��/��YA�HA���b�
� ��O+=����LȞ��-52`�T,n٭f�_tb$��!���}~�����l�LQ���9y��݆fDp� �]:?��}M���Ǒ`1�^[5���\P�bu��Aч��A,�s��7�#N�7G���52|7��<=}S��i4(�D�K]F�\����9�=���YyT�<~)��ft�>�ּ�,0J��y�Zp���@��.��ΉgS��R���:&��C��+���`���"d��*��d`C�'�]\��}`P`���� ��*NA��hj����E܊���ٓ���@
�nm��J��%s�Au&�%WD��3��Z������BB�{��V|H���i[8z�k�	#���w}��]ZW�b��G:�Bݭ�R%��������JB2֑P��~E���P9������\�d�������E�b��)���g;Wq2���6�=$-5��w+^O��R�%�Oi�^��$ϕF�y����:D?Vi@h�bi��o�P"���t��� �n��=9�{�d6fZ������i�o}cԦZ��~@��\��v�����#�%,��x��Ɵ�����9S�O����`�aV�O�tBw���y��Ƞ(q��"����"O"�?�[�p�p�RF��gC3`f��#��F,O�K%4pp�>��y1�)8��
����+��o���غ���8Ko�8V����}�r �J��L��,>3W��Fd�K�E��Mf�Q�R���١��nt���E�"p:(�-9�Rb�M��h,qU�$F����_����%��"��[ӽ�����4k�ղ��%g4Ӓ�tp�Dj�rs��	�aT��T��'4m1����`�+�48c<?���2��`f4#B��kJwhnw�X�[M�!�fsԃv9�k	�ԂA���EV���[=�:���Aiɨ�TdA�N*b!�~
�:�Zu�H�b@���=dZ�EJJ��YDƀ������ᚷ�s��!�g���[w,�f�D*����qU*E7�cAi�����4�=���������Ax��uw�4 &�^�'�Q��]Niu�ƈd\��NS��ɀfo��*��?Z�T��]�r8�OlW�f��̬�_�ޜ7�fP�c��ҧ|^5�?Z��(ˇe`	Nu}�cp�`A�V���7v�ӑ��yi.r��b�\9n'�AV�j�-�\1�n\���J�"�
e��?�����ÿ��#S�)��kdWb"�c�i1��d܄E����.r06��feܯR��V�ǯ�k�����W֥��L�î�[j`����#˘��HJ�����������=!�'��w��5ր� d��׹����U-�&M��\��=P\_�9zijf�-�{��U���(�Ug�mX�v�s�)���q!u��	�l�p�߳uW�8��� J9��ND{I�=���BhJh%�j�m2{�~\�5(rzӎ���PfG�њ/�W{��/@��0$��q�!��n�͞5���CyƏI�������na֤��P��_N`C����=�U01Ћھٮ���ô
��f$�:��P�k��I��Vg��7���E�dQ0����[)�y�z9�A�v�$�j�w���Ǉ�&r�+#����V�G?����'�B)���OQq:�LBr�E}������`K`��1��z<��HPe#����Պ���Qr��g���8x�x�[�Y�4�d�E�`��.���L�c�����ّQ�d7�jN�CL�	)����e������kM#�^@���J,��K���o0�e����wEy ����}�q�������iI�|��h�������2�(�����6O{-@T3q����7��۷yu#~��j�,`4�Y;�m	�cϷ�v�Bm��8���%��%�A���qo������B�@P����vs�B���h.��@�ˎ3�=`)Ӄ�;x�lk��QɅ�OK��I�/����n^L�����ӵ(�ʝ�b�V�*(6n�q��bb"�W08�ޙ�>n�zj��N62����f0_��A���UE���r��W?��y��v��{&}�`b�Y���b.���,����9p�(� q��~�jdl����o�b��BX�1�OE����Y��v���?��Kٷ��P�b��&(&U=��)u_�_��6h�]���4ႀܾ�U�:$�G{���GYNK�q�j��CP�����X��!�k�_�p��"&�N�*����9�n�#�G nq@=��J+x^�$�<8����SD�x�ޝ��@E���0��e͞�v�ev�<�i��ܫ��|��kb��T���xn���^9�Z�����7󀨟D���d�w�Z���\H�US�4곁�!JbC��[z��^7o�;�{�旞O����}��|�<���3Ç��a�P��fo��a1���c��6ҹ޿#�C�,Ȫp���A���h��.��J'G��)B�S
<\nj�¹��k%j�.s��4��5�}�,Ȝ�B���t�F��"?�0�vW?Nf_I�?��m	:�7aU�z)����thI���\7�޾�T��׋��
?��V7�$�z����ɭ�觊�����
}�S������4P�H��+�o^-w��D�!�Q��V��Pߺ�>@�⺖����s�ϰ�e�g�%��'����=�j�ζg��fďsˉzW Y*��1�>$f Dx��{�q᎘�
s�FKk��a�B�F�aO	�G���n���F��>���0gEx\�;�����]���i�[6ˠK�4��8���;H"���~���MP�%OH����M�Cf��o� ��s6��yq&�j�T歫[��^��A�3�KSS�^׆�HgӨ�4ԃl<���y�Gfmχ�=H���&� ��2j���A�X���z+(��͇<�èb�)x=bth��$R]��# io����m*3I����0�NPz�>=��4D{��3���(g��`���!�Q'G��5�W�_��|��	%Q�#���5�n��D��R㮪�t��-E�W��?�M7�C3> �Bn�
Oy�U\�9�ָ�L�Ń�jm�b��)D��.LT���Ί�=G�A!��'f�#�O^��Ԥ������7zҸ����+Ϻ���r��-�Y�"zk�z}>�5�a��3����뤔F/B8*��!�2�H��u�@�iOd6��Տ��߾�MN9
�+?�etJ��4���;��w�/�J$b|�׏:m�C���MyX+_�鮳�-�B��7w��	�J`��\���uw�Q��(�-߷�ک�+n���G�]Q�� �����
�9Tɑ���YY�^kKѸ!��i������6�'R~�
�Vb~��:��fAD �<z|(�z����T�	-���๦��Q��}L�of���T��fmgm��b���3�G�`8.,�=��ż���쳿� ��rŤS]��D&}>�϶�ܗk�R�k���Ee�{�,���Wv����[�6��U��:��wu.ln̯��-�>f�8���^�ػ9z��pJ��Sz��ݍ� ��	<�.����'�Q�����j�E�J�v&ɥmw�A�ef(0FB!�ڜ������u�m��mz��Dڴ)�3�������~s6(��b�*Zp�,�v�3� 6�``���$`���Da�d�2>z��?K�������dI�e�\!&�vʵ~<���3\Àh��t����)���oO��*⎬nO��z}���$��=�]�z8�OU��)�Nأus�!��
:	�=8���u����)����\��`��<��1��r��4R��Z�{����W ��4�^ �������!������	��w�<��v�|�{�
�����鞖sfzz�	�|w�mw�.��wZ=6�� �ջ��h�<r�x�D<n�͸��^�����\����=C&�vs�rȲ�#�[��߫�X�����u�.X�a}<�h(�/�	+%�q��F�֖1�U����	ފ��!T�\I����.`'D�ڶV�s�3��y��i!*���DL�B�#շy��������1d�M/�$�4�8l�{��&O�f�RR��{�z��wf����'�n��k�����������{j�9їӎZI}�S�˳[M������q5E5K�:�A
��sdwǪ_ie%+�W��0�5�"F*믖��և�H���s����_��-�8ǜ�~��`c+@��7��x������B���Z�8�m���j	�wv�q�!�� ���æY����|�1@dc���$�G��t�B�{PCSPɏw���4�BJ��C��җw��r�Ը>�5F�㺫V^>�G�6lY�l��@M�?D��kえ���>:�/I���Y����pp�K&�����w���0̍[We밚��:𮦗���.Α�\�v�� �TZnY �#�]�&eL����H�A���x�x�y��N[��h'�E��V�Zb���-D����|���x��	���\I:Ǚ3��SC��h]u�%�^3�n�u����#A�Y-G¯�s�����Z݁�����5�ߔ C7���$�~�C��!`�42�o<�!�Dvmr�dXP���y+���:��O��RT�Џ��hh5��x�VeKh!߶�o8Hi�Aꕘ�n��.�qfK��K��^��d]�Jt���`;��AO_9�e7M�4�s�Q@&�׽�L���7^��1J����:����%8^ RS��������{a/������W~����#��6���&M���mY۽|ޓF��I��E8���^�e�e���#x����ߴ]}ᐩ��
��#ף�������N�x���0��C�o���!A�M
�m ���]����>u�?:��zD��q�� ��֯]$
�������������ý/�P#�0֜�l���yno��q�8�GE�E1bE���K�D�5u^؈����9I.����P�D�����A�}:�Q�<~��8��l���k����k��J�if6*�Y3���>H�JZL�#kc�������R�F8�0��$]]]u˧@��i~��=w��x2�̃{�K��wM�9�^m�����.��]�y�/犞"}�̍�v4)�"
��.S5�˔O-�&ժ0ҥ5%o4	��9V�CYhw��KC>�Ee�gc΢5N[}���=q,Z�z`"��h:�
�J�ݽ�ܽ&8���:�`#~>ݎ>RQ^�C�A�ʿ��ڬ���5�o�E���fg^caipL�:�7'�Vwvv
h���n9�ӕ������<�~y��4>az
0S�pRo���(�/)�b����m��I�0�L����5T+H��z�>VĚ�$-��kXdו��!rm�T9bZ�������? �{S����+�l}� �tP��Aj�d$�sa̕�&5Q�3�&鶵��3b��|�죘�jS]�7���9eH�,t_��ٷ�J͛[r�QD�����C�lXp(�w񉉉����;��zY���!?��OQn�A%�
��YY��3���dd'�F�괫eddP}	��f�����Dx�C�l_�޴[��b_�2�@�3+A���YCz�?�X�.k�G�?&Y��`D�؟�L���+nٱ*J]�����q��١B6s�/MT�Q]�I��*D��"|e)��%�#�r�WQ;rC-,[؊j��a�<7wwwS�Y�OxH�E��E�$]D�?�c�>L��V��oʗsF��L���zvnH�W�"r���@���<lדwu��/:�����J�ێ	�q����*�^ ��;�+8��/k�̓�j��Rr�]V�$z?��qD�uB)�<?�d� �^SZ��A	'Dnjl݃�ˋJln+"Ȑ+�4c�P6[*#�kf[�q��j��9ǽ�#�$�N��0�*��vP��x�6AH� 9K�	�ώd��xˀ�'�O��,�Hn�~�p:�9dn)7����5��_�2>i����\�d������<����o�7��9@�y���f�T�<VS�8�By�rP��d��ረ�o�UPQ3��B�a�0���͔+�p�ڎ<��+i��zA�YdA-�-ftH���&�*O���T�˖�7�d��O��GJ]��5wx�ЮI�.}�B��Wuy�^81o7|LT��D��ϼ�l�^'ދK�d�`��X�� ��)cy�,��"f��IL�֥�xgAo+�2Ej����[}K�3����T,���W��T���c届�vc(�	���(�햙MS�K9�廻@���~.2c)�����=K>t�>`�q'�d��O���.C��H*OeZ9�>Am�}�y�{X�"Չ�������uC�廂wN*m�JN8@~��X��bE�$�����a�%�
%[t�0 �(@�ӫ�5�U@7�
T�|z_��/��rY�1	1�kq���}�7����������R������ɘ�t3#���٢���ྍ��MT��:�^�a�:�2��"�ܞWu�7��/�3/;h��a��|9�טL��k�$��ׄ�j�R��G��c�~
v��L�Y�t�p�Ƹ�E�۷<} 9��{-���]�L�A���N�d��++�`g�h���X��#�t쵼��du�.P�� �xb�`�S��H�%;�&H�<,��Tds~G�#D�bF��v��ho�R��}�@m''��'��?<� �#�+X%Xg��r�(?;���ճr���jw�V�²O�q�w�MTE˂?UG�(�"h�.��[�����;�N0!}�J�G�,1/��^AbІ���˿�8���a��e�FY�3���;���܃���J��s\�����v|{����n�(-�1x/��V7�l���
��?��@��}��7�����M]Zk�[I{���x/��KvT_s�	���O�1>S��9�*=Ls��>Ϟ��[�EO���_(�v���#�2q�/��}Eh���Po�N��ozJ�+�(|~?%���'�c���~�g�V�o�9�:���#w���O����-�"��sB�5M�j����G�b��w�`"L����[ȶ]5���.Zs�'F���ԅA"5�zUhuϧ��;ᬿեA�9`�ć	-�Ԇ�l��1���.�5�Րy����삭��������L�B )N�7���Wo.e��^���)'=�h�D�k4��s»�c.h-�����ףc���h�H�l�#
��
�~=���1ӈ�_��-N.�zD�7��It����t�cQ�
 �$!eE���:��B��bcʈ�nM�(n �$
��uZ���l^;`�2�{�wez;`>�����]�F~+��_�*E�r^�xF/���\;lx�N�G7�7���I�ȸ���%�U����C��pe��KC��G��3��?
L6�#=�ʶ!������:bh�?��F�	0?gZ>{ĵ�ckK�g�c]",�l~ $��Y�wl�ԾX<�vh߮��5���dh��0A���MS�L\I���׵?R ��&-9@���3�Ƕ5aXvN3՚P?���~/�2/�]���̟�މ��.ӴQ?�v/���H��/GyԌ�r>��VjZ�%��}&����y���X�-|�x���I~��,��mЕI���g6xHxq�a�<Ȋe��n+������1^[�떵���b[k��a #d�����3ɪ�d��X�+灟�,��]�GO�j���\��/8O:���Ž��l��$�r�_)�:����A��>����>oTOM3�Ŷճ`�Xc^m�Uk0=۽9=[)I���w2��a\�O�C?�Cn##��_��c �U�V��Ύ��E�ыv^͏�F��0hq�}��
q�:>��:��,��L��(�^u�[�P�(B`�GW�"��D�7�v�f8�#$F����h��߶	�
jT+
�i����<;V�t�r��ʵ&��y��+��R�|�3����m�3��k6���L�%�C��������T����3&�}��A �7�N�;�8�hԓ�i�P=K��S���?�4����Lc���'D�V���N=���~��4e[�xV�J	2�܄�`�n� ���e�k�?�?sj��.].^k��tğ�v `A�?N=I*��k"��(�1k�SE��R�B�d��9�\d����@�8	�-��q4��	'<m_|c���Z��|�}�}3\�X������ D�i@��a�W'ǚ�od�����A��ALB31+�Is�(�uׂ���CX����� q�GD�bע!j��G�z�J�|gΞ#�T,���'���u6)�EQ!��VB�Y�ߋĪg�O�KQ:!�X15���(oY��FՓ h>�9���]zy�sSɴ�Y�37� `z	�X�)EX͛^ZLN�\Wt�lV��6�}�/:��c���I�w�����:2nL�èȸi��ʷ6A��%����i��e���Y��_���[�u,�'�M�Qr���V�)Wh0�nk�6���&�׋#ߘX�H��жY|��`hB*��j�RFp����d�Y�Ż�"���'����Hg,�7�-��N%yn�S "ol���{o�F�8b]���j=�N��Մ(���[!��|?p�F����Cl�b��@��NBX��B��=M�.A$@�'Y��ķ#O�(�8F��le��`k@�G�V�:?BR|��.�5>����Ӯ�`�;˲c�&?留8|���n�=�k;�Y�=���`Iаk}ۊ����9x)q���_���$��rP�TU�H�/��RO���~đ�z8	� aӁue�ܡA_�r&�g�J��ܣ����"1
LU<�Sۉ�5��˶��,j� ��8�<��{S����Z��Sκ,(!P��兮��b
�FV���Q#� �
,�W�8������v���(����_�������x����p���Z����"��[e�?,��}����_�9�FM� �2�>�T @�1��a�Ι�=�π���(��@��8��	#��A��P�p�|(�����sA��|��S�� .2��OV�s����P���
�>�P1W]����?Γ���l���U����cX�U�C���J%6L��3���a�f}W���;�&�`:��]�eYX��ri%i��>;m�8��vM�T�����2<�����<�暿���3c����M��H�<��@�&�}�\�ĭI8N�����D>�A��S��PA���I\���6m
s�gO;���z�h?>�KCJ^���\w�L=���\����Q�{��؟f�t�;� ��(���\��~k} �kM��ٸsQЖ������p7�*��9J�y��[������
P���Qf��Q>��ki��R��1�h�d���"Ku4�[�5����G ���Mc��ŋ1^�x�&7��,�DwNFF�y+_Hf�%Ƣ��[��q�j�����V-�Y��;�1'ry�?6�x�����&�Wҩ�"#�Ĝ���
�T�U�Ek��ï�'�������ul�_G������D�0ṕkD7]����_������3�Y#x���Ċ��d_������*���!�X�_���aZ<�8�Y����9&V�9�Kz����VW�O���z�kj��ϿԂ���m$�޺?D,����f�{�uۜh�P�}ݼ�╨N��>�RWjK�n^i�w�YW�H�'�	�\��i��"4���`����N&�e*A��B� 2'%�L���:��_�����s����1)�+�_~�nl5��|D�7�^�E��p�4]W�`EGm���eԑ�{�f��Wt�f?!{��>ߗPi��h��q��fX��v��v��j��e�)�w@��S�O~p��m�b$�+�i�>��%. �@�2Ղ�=���A���v�vK�"��&��Z���$�2�:ؘ�*ĬK-��Q��[7�#N���>���Q.4��q��]��ޢ�!�����Kf�l��p�o��0�,�� �E��v��/��}%�Vޏ�ȃ[Q��_��PUb?�s�g�\���e��.$�?BX�1?�m�|]"�3!�R0�TR��K�iBC�eHX_f_j!�!�J�l`��8���L����Gs���qc�oxQ֬�N��\�y���Nx�j�`��r+p�fj�t��H��$�zPGA�T�8��;���Z�B���}㤬3	K�n�#�ݮ�X�l�MC&��������H	�����}�+q/�Hx���-q���Ce<+�X��2�����n�&Ѣ6G��2�5�ח7k�9��C�ͩ����ɐ��/����*��Yh�۽�o4Kh�"1B���7�LGp?���z?o6���ح�И���q���F�dxm���`3��q�Z�R�:����"����~{Du�[#�P�#2?{�_�*��AnѶMxS�H"�Z�B��C�&�?��S�b5�D���>���WQW�[uLXiC�������<Ն-O	$��/F�՟P|�kA��e
Ҹ�M��]����x橆b�T��C���021:���-�����Ao2jc�
�`bR~`X��+N�N���H|*�@�o�ݜw�:2:�vlV��d��l�k�@=!f�G26I�QX�/Jra�����{6�4QF���^�����G>W"G0zs�qn|�t�C"�/"�1ˁ�`6y��6�����.,��[#�Z��D�����>��5UQ�ذ��-e���l[+S^�|���A\bLπ�P����S�O�5��Rrz�_6's?���jAp~�é���cC��7Y�mCU
�Gd|٬�/~O��ي�D��aˋ����CH����J=������W5�E�f8����n�ѱ������)���ֲ�w��*�A��'qQ�w�����R�x�h��#?�~�7n�����ٺn
4=&(�̓T��O�!NnRh�ciƀ��X��ÃKP�h��Ԃ�Ǆ��"�<A-�DФ���g1���%b�1D��i�����b�[���)~ݸ��	 ��o���R%��اv��?��s�����]dJ���g0�y�/�>�R�&'���c]�+���fx��j�����2�pq��q��%贪}Ra��H�ӿ���S/��[#j1'N���`Ǿ�:<L{8

�>$�����fzW�p�:x����8��\"�Xbo�%E�/�qz)�-[�Gp����6����FeR�ì����Z����'�YK\1��n
�����͜"|���p�p�=˫��~�Xz}Q&�	�m�dx��hL}zq��3{��빞:fPy��h�U��y�ӛ�i��W�!�b<�.{J�Uٜo'��(ة@��)�(�i�i)Χ�z)�zb�3�5��D=1����n��>�/��j�����f����M"Rg����	��Fi���d� � ��L�����SM%�61a���e��]�%=�ɱU����?!��Z_N.P6~=�u��^�o�X�U��%����M�k~�/K��@����r�S�+�����g�v.�z?bQ���q��u�f���b��a�����ݽ��xi�n��Z4�Rmw��.���X��o�ˢ�kM~�_�9+����o;%i�f�Gx���x����*��酢��	b�v�s��k�[���9uگ�v�[���&"��}>�+�?��bV�cE��ψ8��ao�D�szl�V�T�:�k��o-%Ġ�1I��rc�����آ��bKaM�Ye�R\�kM��u9��1+6������p����~ar�b��U3�=�~�䓬�esΝ��{{w����T�Ǧϰ�}EJ�b���'�[Q�σ[ҵ��M�4�l��߶9��	֪6�p�x/.3g� ���_2k߸��o�k;A��P�C;+����KOn���'/���mcN�T���4��t���!'L�L��6�R>�E*w��s%�|�7��[v���{J��_{�XX,����f6]��G��o���Y�m��5i�D��LG�i�&6	`X�	�B.����]��y���)�xz��ܶ־���rͬ�7w�M�'f|�Bz&ȹ�(F��¾�)6������E�ej�J�����g�������;b}a B��:��\���?�ɼK�&XoBj�g���C��]P���H�G����ǁK6U$�\�
	/�����3���a|m��B�Z�]��:����c&&�X�+��NOd澇.t?�u�R�<����j)PH�Tϲ�$��a��t��<��� ˿�d�� $ZM J(*[�
�9H�Ge���@J�M�Fm�X}k��=x��k�����F�'�cg
�1yR
�����"W6qg�� ��a��.�T1s2x�����A;�'��h�C��ɬԴm�*�B� �2C;��ѶL]�Ƿ�!����X��C����d->~G1�F���/�@�����}�Ot�����dj�1:��@�4�X���Չ��{bJR�D=�	��Ʊs�C�+��׵d~���<u@\ө�q:��s�xn�0���^g bs��}�d)�,X�t}����o0�����k1�W��k�[�6��0�V|^����7��2�����l�_�F�]�/0B<Zǜ�S�/ �!��5�`q����o#m��c���-^�j�r��-3<� �����U��88��r����ڱ�m�n���ffOA{�Ԅ���p�>������@p�S�X�T�&�*	�vZ�&&ވ�3y�4<���[f�eW��������&����^����X����d��;ʰ�� ;ݠ���� ��c�����;���rL_�G����6& p��:S�d�_��<��e�MH�~<f6~Q`����f'�ʳ��Cý
����4e��aT�v��*i�p���NB��ޠ��@N����h)�!s5�:�1���*o��i�%���uS��W`ʨՊ������j�G ��sF�I����we�$��d�!�Z4�G �=��HB�+\<�진f�Ob�����y�@\pMr��0ˢ*�#A\�#�^�3�D<�pkY�b����PW|l�=� @e)�~���qG�;��m�'��p��_��ݧ�����gfwd�Ε")��yj/z�l�k�,ܕhň���=�5���C�2m_K"f�ըR�f\��<�C�Lb:u����I�q�������������@'O�/{+�᮸S�Z��F��u
�b���g��� ��r�Yq�[Mr�J�{^��7�h���]���C̬��V+'�ׇ���I�����m=����n|�#*���C�x���"�ȆU�����
O�v%����4�����M����f��t`*v,"B�Z��NF�̮Q+���i
��fH��rǫo�p1E�[���k�$ΫoY���Q��o���Dh94kR�s�~���K ��G��x�t����J�(}G	�?v
r�^�d�/�lа��`+�$��Q�U��xm�y	$,�H| �yz;@;p����^xI��a�_��^s�_�D�{X��^�1+�[��0PO�>�ep0�;�S�I�e�o���^vj\�RŬno��_p+=��aT�7i���ҩPt8�9h���`�FW�R��,0�9���wn �é�����-Ŏ��P�1�v�[����C��)^����:z�'�_�dH�V��l����^�K*��S�z`�ṙ��8�PQ��	�A`��3{<�(����������v���l��>U�����>L>�sG�.�{�4�V�z��V�;M�
|�§͸��r��K�/��o���M�ד�U��N�����po�_�����4���.���?mR�-^�fױ(����Bk��u>��D,���?�
bY]��F,z�Q⢎��B��D�F���q1�ΣM��+�\h���B����"�ܣ��X�q���oL�.Iܨŗ��ŻS|�7�!�(�g� ��)�I5�ڦ�O��H�X���Zq�u�qA�Q���0Z�
& ��q_j�J뗇�~�AI�a����IY'�"�5a����n�Ϥ������b��~��tCwȞ2�:��S��S��_i�i���@�Jߍ���Y!h��N�7������Y��
���$u+���@�w~W���AT��6S/c���l�"X�Y������R�^�������q�}��&����Uw!:~3���R��B�O*m�'�_�I�Y�Ib�_�T��F����X��@:���O�L�� T~�s�Sw�q1��b��YT��"ԃ��r*�s�)��n�5Cq+V�,����N@I?F<9�lҹ�����t����aJe�D]������|2Uo)sYO�A ��������� F�y�I�I��^"��Ľf���m1 ���q��S�%EUOZGZ��F�;�jkpωP�%`I�M<�	hjy����#ǉş�@m�}���쨊��/��>{�.�/&�7�Ԛ;o�$��� ��,E�T��k~� O`x��J}�f%�����;z�Ol(�j�t�2�|I�} �d4)4մ4�;Q�
I�3��9}'n:aXex]g�d�mNT�qx�����;/eV*�Y��� S���+�C:<�V���.@��Й����������8���W1a���q����_}~��`��>|�6��׎U���FGY�1O��h�VwT݇��ȅ^�b��o�d#Z���0�휳E+�� q� i�C��}���p7/<��]{�+3�F�ȼrG���s'������&��jAH{�߶�G�\2����0�3R|(�b��TsJ��5�Es�c��ir���r�:/�m�y�J�mS�jJ�|c���F�ޚ�xV���;)vE�f�8J�*o_��پ�s�1�)�[͍�DK8��<�*�H<y���W�c����<+�	��a��� 3J��S�(v;��)��I�rL�&�����U�)DT;�%C�%�7��j�����%��9����r�P�e��b+�j�����}x~�șH�&�AK�MP�u�N3tk��R3Y�Y��~��=3.��?c�$Un����������~c�A�qw����F�h*���.]�������z�;���|�P�P������I>]1ӣ���t]J�$K����ᓑ�%*��f�-k�f��H�0-�':Wlf��]+!��u4����ڻ>5�ae�����F�<�͜L��1�o�,��.;��S�~��3�<僦����@����Ly��w*�����Q)2"d�y>��4apG4:
��O���F�� )q�0�̄a,�,��ͦ<�?�A󉟑Dp������oĸ�gLA�>Ȥ�Fl�X���{{J���^��afe��]�	j��l��E��>E����h�ڠ"S��u!���s�*��*��LZ4S��O���݃F�pp�:R��B�E�{�*L|�lQ�}:S��0�{ǂ1����$ XF���ђ$��`�e,ś�Q-�b�bn���S�cFDʼ��ĐE�	��x��wX7`|�����~������Y���Y���i?'����K*O�澕~8᢮��h_�I�h��8>y����e�a��q�.���%ts䅚�VִTb.����v�e�(PbL���^+���[��s4j~N���)����Uś�����x�F�������o'�������[��|%��N4c!������p�0.��ɳT5� �Tb���Ý�'^�A	!Oq����S���鏓V�
܀s���V��D8�P��-�}�����\Չ|�O	P7�g^�_}�a����,��w�E���i��"ˋ����/*�����$���L鄅���#��nm��b�yIb���L��E�������Spmƻ.����5�$��Rb��iA��c������
�Qtw��ʇ���RP��@q�	K_����K�յ�b��H�S솖�̀���N�=:�0D?�.���(V廜����ʁ�a'�j=�1\�j�$�@�l�Q�ݙغ9�lh���l�U�V-�����9���w����/�3���ܰ�!�O	i��a�HE��_��u�#�-E=�����D+���e|�Fw���R�,� C)͡|�X�ǹ��V�zʂ�`����D�퓦:�+hӬ1�����?��E��K͌�W��R�@1�R� �{k��ܼ� �KS-�����Ȥĉ��uZ��1�1�E�
$-�]����ϥ��V�	��1�V��{�JU\��ˑSM��9?�lsw:���6�Z�%�W���	���q�Po=L��ݼw������\']Wq��/��@�%��\�3F�l���$��pHQD���m#��Z;L�n���}/o�}؋�8�ˡ!I��l0�DSuv�\Ϯ�Q(��/���*:��]?B��|���	x|�ꉋ�)���-�|噍�f	�����T�E=�Y���;���3|�v����õ:�R�]7)��y�k�F���1�@K3{%��'2+�0�����~鏏�=�,�&�qkm�Xy���*�r��w$Y�3�������J��]�zFX��?i����a8�X7}yg��ϐ�%L[Yͧ��ˠ@L(1�]R8�}����P8֋��<�7K�����B=	���{��!�ԾD	�ɼǖ����LB2J2���ƻ��:�'�6�;�@-�ncw��♩D� Ӑsʪ��R�:�bCT�Rӛl^��X?��O�U�7�+�x��Y�Î����=S���:�'L���� e��=D�T����s�XT�c2]�]������@V۲͸`�o�U�&�eOy_�D��J"�	4�YaB/�ހ����0el���x�#@���԰�ЃfZv�LS�}�p�	���@ؗ���"t��� �;3Pu{�F#���;��1>���X��@P>N�"��ў�8��&�3�Ej�^�q/��v�پ�gED3�3c%��� p���7Z���o:��	M�m�单��p6ٗ�m������Ð\F�F�-U<e�	�L�{������1����M��;�II� s@����W�g�f��@����'6����qǹ-^}������(q�	�j�P}���̥M�� a�����[ݰ�6�i�ڢ�ƍ~��|�H�޻?�m����.x�Cѵ!og��;]�,
�]���My��Pd���#��Xz��/F��
/�֕��B����^�bcK���&����M�5�4ԩ�*T	��ʼ5no�R^��Z�.��|R��%<^�`>��]U�����P�8�e0J�٦s%��{�t�\��f��J��8��d$*Yu�8��I�%�����6���=X�o
��{�
H���*���)~"&������+z��61�&S(��N�k�b2�k�����
=�*����\̓�v��>�X�y��WrK�f����{��Qq� >��{m�⸆�(�_��ɪ��M�$�aDi£��7<�IZ/��;��\������IAc���L����0ӹ}H�]������|~�Q�M���n�s�y5��N�U�HV��yW�Y�#ݼ��FZ�Q�a�bGd�un���,���I;�X�����0C�&��O���<-E��V�$��
�j�"D�Z�X{,i3��7MS2����C'L����"��Jj�q��8���)*���e�BQ���+s`�/�X2��S*�s����d5nO�-j�Ck��f��$�lE�I��� ��b���S�zE1 _�:�V�����n��#�S6�"
��5)仴Hu�5�~�9���������X��9�+}!vXr,�n�!��N��!��en�����S�l��~��\W+b�?_q��+ܮB9z�X�k���W��I6�v����{��g��Չ���r6�wv���@aũ���8�>G��Ƴ�
��sGs�ѓɜ2�/��G_��E-�?]��4Q;©x	����1�7��80|�%ůg��tbk�?rp�\x={�3+.�Hf�b�4��Qv/{]&�MK�	��r cq(I�9�>��x�J�`!�+u�"�"&����
/�mKkZL42"e��e�,ģB����מ�v����Pߗr���+�~�е��I�w[g�����T3���L�	��<�o�����}gͳc&��R��Ϸw��Z-\���{	���Y�u26q\�^7bBg��E�O�V�)������p�΃����k{j��|�N*N/�+�%��ϓfח;��{m���D5p-�EB�L�j��.{��[�4�M�l܁meĀ}��"b����s�N_�/�_m����a*S�2K�q�/�����R��=�9$�l>9�P]K |-�+S��U4.�1�g�,��-df�]>&�%�{>�W��&Q}@1Y�"�p�S��S��/50P�q�j)�ٍq�w��p��ǚ�#��%�s½��.gҫ-�u�T2ř�窩�,h��ؗ�v�����d��+��}-B	��_-����d䌉��l����\�2�GD��_���Zo7LF�*U+��%3����@�Q~I�(�֤2,����[�����=�U�+k�֗��!Ƅ��"W���"��w�a���5����ӫ�>�b�x���E���>���@J�%���U��	S$��s����:^P']#�<e+�H(��3��Si��DE�Gdo%�����2"i�U3+���.b*��K�bˈ��x[�$�!��U�a�9�����O�V�A����@Zr�Y_���zY}�� pp*Qqm�5WdEO��j�H,�{���+�����u��&Vr��v��倭6j
����$=�,��P�s�7 <�Ѱ[ھStc������Ƀ2"J��9b9d�� 
��%�х�
S���۞Vآk�r�r�������0bt|ȗ?rZi#�_����!�7rW�LZ��ap0���#��=�h���qS&8�r���ۈ^��gOr�	=�g� ��٘�,mƚ�Ke����0g��b���V�4B'xl�-:�Ob%f>�C�+]ƅ��R�ˀ���~��i����v����.13��s��i
�����u�{�Օ��_F;F��4�5Ƚ�&YV�ѻ̕oґ��ں�ѯl�+���'�]�o8��`����f�M��$�٪q�o���C_k��-�o���u�W��R��\*߻�%��!����網�*�!w�]W�	��|(Q$�k��Ŋ��w���e��ŕ�	2đrAz�$.!8>�yN��q��>���]L�:�u^�������:Ԧj\A&�9ьɠu�
�-׮U�{�UG�*ꃶ�D�ĩ��Bެ9��<�2q7�qm�V~���m"�΅q竔	#���H�[z���'�?�
�~�����Vp���8��+�N����T� _v�4J7��qJ�"m�#�B�u�)Ĩ����]�>�^tL>H]I�m�Z�C��ί3��|H�@� ������LZiy4x�l���h�/`UV���.��>�%�ƗY��2�oܬN�o�(\������p���8׽.'�b85S7		�0�L(Fq;&�Ti���C�X��Lj�\�G|��
@�������$��&��������!W��W�q���CD������!���S؄�� �!oM�0��_�qBԑ*�0��+��q��7w���+I0Y���.#��|�KW>O(4���*��l��$`F
?~YP����X���4�t|�@Y&��h���3g��������[d]�ۄ��-�wsZ!�9����<�鬚�,�$�ۭ���8�O��l4ix%f�E�ۢ\0��p�p���
�H�ĺ��n6��D�W7E!�PBJ�����{Teg���K*_=��?t���5�<g_�L&r=m���=���r�On����͗S) iPW%3�#!���/� �z8�}��T�Hu
-��4<��?���o�$�O��U�2j:�)�Y���f�>��*p�)y�HPݮ���oF�|�n���es`�8�ʡw��sWy��a�؎�� �q�ƹ�`��
5D+F�Y6r�N7ui������ʛrxCx����u6u�`�Ii��z7�F?&s�7��Ӹ�n��`@;C��D+'/���K�'z�+5�����@�R�S!2+���v� "egD�ՀC�{No��^�y�	�Idf�hU^��z��S�H�8,1M�%ͯVbO^i�%C�O���2���|]Zo�r�ϱ��R^����M��3%�7p���JƎ�:P����mO����v`P���	���9F/=%�_n��~�䪡͊�1/-V�I����Z����gw��	���˔��P�s[y�S2zç�*�����X�j��9��ӌ�jI��(g^f��>�/�|1ė�{�����7����O����T�d=�=�w��ã+�]$lZ���2����2��g_�BȉE3���{wt!D����d��������.l�!^�s��u�9�b4z�kmZv� �w�- ��6>��;<�`�VDX�|ΌX��|AoJ}V��T�X��ۧ����)��C4��!�;�C���h��j=�44<LU$>�8�O�ܛkBC�|oy,�s_�G״������K��!��]�8,��	 ������]ߒ�y��W5S;Us�̱���9ݽL*F8u
R�c�.H.�h���Y`��=2"���W�,hh�������Z ��BM�-�q���ԡ��<�������ۋ�ݬ`R�o�`���7X�4ނ*�S�`��R;cQ�mB���H��h�{-y�y� 3����jB�]07�)60����%m/BхСTc�ԛ��6�:$�g�|[�Bn�R耠H���:��88�?��i�!�c�ޞ�B�?Z��Ю�A��6X�nˡ,��6�_����&q��󰊂���!��}yC�=F��.-i�#˩��|4G�����0��yRi�?t&妇��:x%O��q&t�i���u�I��i��*T�4��z.7K.�	����Va"�lj�Aɢ0���� bH�Z��h��f5~of~��8�@C���!�N�J�n��Ӻ�w�.~�v��5/���.:�Ա1�Z�+ڠ�?`S�� �v�Cݗ��E:��,�mt-m�R�y"K*���������l�'42����![���T��*�.&�Z����J����������w��b�?���m/m��q��@Y��+��n���'��e'��<��nW�K�Xc�CK��S��}B���.[>�q��gFk�W��#�!#1�ٚC��q�>�;ҽ�Y�ج�E�����2k.>=H��2
vb��*�>7�%��2�	��2@o��fG��7�//%�yGW
r�jW���~T��Jnxoxd0�A�(_�,���ݧ�j����z�ؾEA������h�][��w4 ��}�,��mM���no����ͺ�� ���ď���c�cK�L�w;�ʆ�A�՟���vSʄ8�Z��s��w�]��>.>;b��U��v��n`��-�zac/QJ�|�1��E>Ԗeu��%���=�."Jun=,U���[B��U繺�έ}\��_�l��n�d�u�(�8�5aپ^�ͤ�W8�e�Ü5�G����$'R��Ow��u>��ñ�z��ng��k�g��<�T���}HWpu�wJ$���:q��tBe�]v�9W� У�}-l���Gcُ ��H�������[���9�X亝�����u��V�Zy�
��	P�^�l��RB:�BuF�� ᕆ�H����~����ʞ��p�-Q��M��'H�)���d.�s~���?�R`���>���Q�@o��x�`E}P�.�iu�ab�+&3������݄z㢪��qX�F��!��Q��;��4�O��Tߙ�M���=r�O��)l���~� �.s/�?��ݓ��G���r��x�7��`�شc�_�M�i%�d˄i��:\2s�� $��sڎη����B�����<��I�����W�/����v��6����.1�:'N�1�Vڷ!�o�b��͆5���� a<E��S0[�&x~P5V��Q��غ�zO�zN�TE�qcVݯca���f�Zb�(�)�a��&�]���V1lVg)�W����V����aVcT�5U�ֺ��6�E�F�F���2E�HJ��IWx
3aT���ڞ�fvQS����3/����u<kH�x,��e׮�x�T$��Fu�j��Q�lȘoW��R�%�s��`�VyH�>%M���I�WD`ty��]E k*G��%q׼e��T���Shw����av�8�>h۽R=��^��H�~�2�B�b��a˽�?ˍ?k����@�O��\�m"�p�oz����=)4(L}���[�5�gmm�h�Ehr���l��> �M�s�����h���d��!����I�P���f�B4)g_s�����H7!��E]�b�O8<?3xM��]_<3���	#����h�,Nk6]5'0�MzU�����/'����},�˧��O�D1Vw��͵�G��8��)#�Ѳ; �5�� ���^�'����"��%�o~&��լ��yyEmA#e*�1��h����|�B�{`eM�J*Y/F���tis~*_
�J�~�l&���=��Q̂��
�[����Q�u�(cL�{'���$�wġ���n�.� �2�pZ	��Y�P�r����N����-�*�\��d�/q��om(��F��J��/�Nz�=�-YtT4��?L�`&Ҙ1Z�o�N�n��:dr�������2�)���5�&f�N�2�� �*e`c)���AY'����A��Nt�R-�_{	i����X6_��G����,`�3�[�c?��SF�}�Sà@���&���PF"g����޳�ͺc# V�ި.�?m���8�ڦFed8>'H�]�]^��D%ㄏ.��բ�rK�|�`�g��e��9r��ӑ��2��C.��XS���Bb)�f&����8L$4�$B��O��S������s$6��N+%k
m�+/����:Ӱ�*- Ã�x�q�pZ�4q*��;�M���ۭlTCL��D'�r�7�9<3�}O�C���ዖ�9O��:]�k	�Vj���m��� &'��wsW�"���Z��R�.����]����ިU7_S��l5��7Z�'ⓛ�!���}���C��?�Iz��?v �#l���beܐ��p���)hoO!�l��7л��E2c��w��=عe�
���=�C�`�s��dl��=�ҷ0Pt�^b��>�"f|u�69�Ÿ}�(l���?��K������HN��;��[�׊�Q����yB}���ˍ/�;t+��4��|L6o%���,���S\��v�!��I���Ēb.ø!��*�O�ڹ�E5���-.[ٌ��ܼ���蜮?�]�>�5�(��EY��X�l%���x|6�X�c���|���T&�0M}@����7��6�R.���6u$UZ��d�7Ok!�w��2��5��E�##m�Z� ���FkK y�]O7���E�Ո�@�B��:�]tR�@]�6�"҃C���$����`-��yj�ɿm����~ݛ��������hi�a�2�T_�^��Y�������䯂t�顷AA5I[�mb����� ����� �	~��'z�X-̺�n���N-)ٚ/�A�s�������?��q6tp����($t�ǲ��&���eN!P�6�M���xO@�8�$qd�����`h�o
LڜϮD��3+�b�����w;�f���3���ċdݢ��R?��K>�&nG���b�*l��Yi���Zj�龾p8�����7��I|�����*��J)/�B�F_��{��2M��v}�H�@�
�iir�<��h�<��AT�K�x�-g:z���Rtx"�5��
~>�vnco_�5&����xDs/��$h���F\�΅y������5!�6X6�>5�(
�/����u��҉	E���~�rB>"!���E9����G+L�f�KDII�Ҝ�g��q�o0��*?u=翆�H��[��V?�I��s��u���?Rq��&�J)��H���T�-�8.eo]t7���9|sbb�L)�����'�N|�e�M����؎����K��D�a��<m�L|�)瘈!�+_U=�@�QѴ�"P��q�;u-{�_�u���m��h�[��eR������U��a��L�u�p�/3I��3le��RFZ��rR�4q7�c?���w�8T�˵L�~�@�������5l>�&]��|U�-k�ou�On]%Dm�c#�^�u�>�4��i�p�����Z�#�]���$_`h�J�ց�_�q|a���������p�<�<H��eC]��xdW.�3G9�èŌK��8eO��>i%�+��q��Ѳ*��8��9��%���`���{Qݙ��f\�T����1^���>m��h=�J����b�y ��s3�į���>���αw�q�d�)��-|�A�d�e=s���SZb������Mt_�H� 1j�{�����յ�Н�Я`qMD�}+����d�d�^1�@����������|�q�u����V�S䨼�;��&�,��?~4Q��_g�q@y&zb�L�Y�<���g���#GuE��������i�	�*S�����٨)(�wz��'nB'w]�n��$��5��	�0��‍0��O�����1s�?-P�>�.E��E�XqNL�=�'/㍵�qW�qt���Q����a�������$�3�4�ټu)����b%l�K�+V޾�&�g�6n]ַ�ӳ�1��U�����qE���?���������@��(����u����2�'cvZ9�/�R7���*�f���"JI�����#>];�/�>�o���^q�)D�J����mO��/K?�^�i��4"���d����u�Ҡ���--�NE����[Y�,��{a5��V?�p��]�eV�������M=�o�L0����+~�O�z�5Y���\��"�������ֶ���3_�g��qi<���gC�v�s�$�qM���3�T���R)��J&��w	�G�`�7����R<��N��ݤ#;ɪ�&��j<lB���Ƚ�	H��y��|"�t�qh8NHA}#ϙ�Z/Q5�{6Y��Aިǫ7Y�l�H��:��d����K
I� s}+w�4#���"��c�*>>�G��}n��`���"��A��B:���PO�H��)��M0� cQm��X�v���5�N���Ȝ��H!k�2�vr�A��ϊ�?�\~�ow���W�pD:�}��p���u=ꍇ�h���TAA�$��P}oR�յ���^�,�����
`��������s�Ը����ټ��!M�}q�����[xAG�Z���s �V�/�˗�?{�}s�'fOSTm�%���jeJ���
p����	N,�����ʛSaХӉ�@D���(���SE�{�R�˹��7cb;�`.�_��Eڕ��B�����ҽV�{���Zw-��;��Ƶ�F�v�ݟ&|��֕��(T�J(�&,B�d2�H���eJ���6PR��1���^���H��Mt9R馀�G�WqұS����yr�Y�@�x�c�G�<�+� �P\T���7G����B��<qC��}�~ۍ-$����_;�\��Y��>�J!�B��h�ge��Tj��o����+ϒ���K���sOA�M��b�߇� �i��x�
�	����X��
3NA��XC�"�ˊl�z��W>�@����J�R�`��㟁��z��T<ҷ@��v�bM#�s�	^q�FA�ߘ?x����6���ո�͢�1<�d���|���'z�ۤ++�����~������� (�+�r�~�T:�X�tc�R��ݫ`M�]�ao�-ɵ�)�&jO�W`�֞�!0��v�(��kWCJ���M�����W��f�Y�uw�R�5��нs�^�Q�{�X^-y��1c$�?�ר�E�a!$0��q�Y���A=.�����G2*��5���ټr�D{|=h��v"�&��_g{��׏x��jF`��>c��8�ς�d�{���_oC���u�U���s�`!^Ǣ�b�������r�P�컑�߶�&cG綥hyT�m`\+�_����kj����Gb�䭭=RAj�h�?u���	������s�:Y��\J9�n�L��q2����Ao����_��}�����Z�)�iU���` a�����_�S��k�^ƪ�Jf>��6yN=��5l�@{w���Bli���3�q$Ė�	壡��k��x�����e~�~�Wji.r��`��f5V��O�� OO��Fw�~�P��'6T�5`C���x������~�*0va�౛bjL`) rXJ�T�ᬬ�=X��0Y��R��b��B�c�h8�35���w~H���<"���2,�����LQs��W/s����� Q��¼�"�y	Jh'�:�}F@���)�}ʫ���Z���-X5�vm	+��"k��eVO��w`�'M���栁����|�X{�o�t�0g*ѵ�����/ �M�V��@�T3ʱ"W�N/d`N}��)S�K�{��E����e
����Xg,P'e�#���u��K�$�,뫤�?�����D�Z���|�|D+�,K׻F�%�Q�.+C�8��	�#�+8݈�v�P2x��~t��"�đ,릣:E2���)H�1�"`#Ĺ�U�u!��}��=�,;B��H���?͘�Ș�x�D@޹��k��G�c�۸V_��d��`p>��sX�����eLK/�kˑ1;�Lۯn��:g^-�����ﱦ8��F�4���\ �����?w�D6�w_\�1�pk��K~��'��t_��\&X�n�:	�x�b5�b�~�Fx�V6a҉���������d�� ?�FvU��x+d���H�f���&�_g��/v
���TkX��[F�z��!iu�}�*f"���6��{~���ȓQƧ4���a|!�o�E]2U�+.����+W�|��/�٥�yi�1�>��ނ�$�?�ῄY�G� �Gb�����6G%\�ޔ�k�OX�[�m}��p{�+I�����"�^'$;xl��%a�h�#0�X�I|�/��]�G��A١��(Q���-eEBm8�-��|o����2@��|�.�ɠ������T,h�18#��\�9Az�x�N�4�Ě�[�;2����}b<x� /��^���i�M�>��2�ȶ����6�)�e���ɯΝ=N��%��{���Z���NT�d��6������@�z�E'Wo�ъ�A��3�y�a��	�E�Of�Ѐ��� �����Ȅ�ٸ�P��^Gb�$��Yj�W�ҷ؅j����k��U��د�g��3C��G�A(�~9�^��Z�6����I���o�)>[��3�gr4c�@��je[�;�©���?�ى���p��IR3z�-{���R}�ۻ��م���vfMg�z��ގyP�os޺��o����?i�F��|v� �E�@w=y���zR1�S��t�J�6�0=%]`�N�;a�0J�c�+�����=)�?őw�I�>���0����$���Y����r�-�i(��{^mla��я��o^n>����&�U�`��h��ݶl��*݇lj%�(f�����#B�ѡ�d 澿}���S���6k�r��=�v�L�	 <+�M���J�m�:��FO�u-�II�߿��voc��MY�O����cIN1�t��0���I�\@gό;��O����c
�����1�D�J�Z�
�H1���_[��W8w\)&|ϳV������}<���.LP����=�Czc�`L]ب���%U��r���~Z� ��qC�]	Ɏ�>8⻞�[�"���-���F��x���	B'���e�am>1r:���k#���?�'�q��o(��q��w��^O��$��~Π�Y�72�d� ��`�=��U��γ!�N�E�N�F9�����"p�޼�(�C������e�؂Di�l>�xi�A� �.w~�z�`bG��OD���r��{�`x]��{�4Q@�sJ���΂���Xq,T���1�FĬf�o$�Ԩ�>FI�o�n���Ƈ�.�τ]�����ƌ&��]�E�iu�c)�ij�N�oJ.*$�EK��ju��e|�ؒ{��'��~��������co�p7�A�XA���������Ĵ��s�G+�/mth��g�w
>���I��>��)��J��wbqb9�")1�K�R����2>`��H �l&�h�u�(��R�B�P�4��@/�Z���AS1۝�?LPU���*4�b��wQ��y{C.�oc�-��dH<[�rP��hF���F?��	X�9*��>�RP:f�e�z�T�Mn�����#ҥ������T��f��}���oAt��qף�@bb_��$Օ�	Ĳz�u�&`ėח��7�D6��!�����W���oo����_=�ll]�F��m��ӆx8��^�����v�UQ�� ���I�_���	��U,���K)¿��m��2��5��y��@ܽZ��F�:"��s
%n�NQ]���\��2�X� X����ý��n�K��f4щƿ�f��U�����Ņ�iLN3��i����ڏl�r���	�h�[x^cH��JL��^�h�����t�d2�nJ!��TwK*t�7�����9Z!�P(�Zǲ˦A���3�W��s�i
w��5�N�ǟg�� c�Q5ǂj���KmgΓ�_~��9�����#m�[�%� ���G`b�u�����/XҜsޮ��b��+�xB&��B��J��C�2kٲG/G�&���q�4�`q^\d80�wA� 7�0Wۉm��N�g��oA&v��?[a=~:���Y���L?hY�T�V�'Ö�T��W�"�۲J�@J�IRd-��u�Z������$�PIT(����HV,A �ܩ�Q)�2�!�J#��Tڟ`��Quxh �(��LO�s)݋�?�OA>��۴�K��0��b�T�Ϲ"hM�(�q����O��pXC��A@�3�y�/���_�{���S��I�ZA�O
����"@z@��SS;��&G���'�U��*z"y�_V�X��ڌ+��T���k%9ϓ)8(4��S	��5&�� �N2��?��?0�8K��g}��,��HM�M���P<�쮵�zG����vG������64�!�.ۓyr�r���Z�W�P��?����7�Q`�/p����%��S��+���+�?��$��#|�򯰜$��������t��V�i�е�$_=X�^���S�D�L��H׎K��Տ����;b;���^� ��>�_��~z���!2�̝���G/�y��:|� �Gw[��<�M��h�4��Y����,c_���YȮ+�ꌢ����L�l 믬'�����Nr
�֍��k4?/���P�dhw?uj}Y��M��"�_�r?Ee.N��L�=?T�^��v�r#��8��=�=~$�a��S61�et�$O��_r���y]�ڀy��o����ﰩS�/|��Ĩ��Z]v���}-=�a�t
�5ձ���ԵxY�vl��.�_�����[4�V0f��v�8��֟����/'#�~L���Tf�G�{�ec�!P8�Q�����Y���B��O��,pE�����"�N壊6��65�$6{�~�2�l���c>�4^��(¢�_��+����ާ!\�d(�u�Yʃ��Ť�r%&P���� �zȰ?��َ\�uϴ﷝�� EsJlQ˷���/o��5'����P��6=��2ZrT��>�8Y��x� Ɠ_��e&�'�/2����,d����̝d`5����a��n)�ї��-��،g��P���k.+(P���?5qn�~�dc�N�].Gc�c����T�L�������%�\��
�T6m����arC9��\:P��.z{��s�tp �����	
u�ϵ����d8�� ?�K��b����9�w�]
�
�8��'7�a��C(L��8��,�u����f �T�9m�]?;d�F�&�4'��cf�_$)N��-��d���l#jat~�j.�JןM\�~�����/��1�� ��b3�8�T$a|)s��:쇅�DD�Xb���?���L4sAh�*?�����>Pm&\�����ϐf:VM�G��22T��rը@�M A*պҝԕ�6;�'��+��T Z2���-Ѓ_�Z���������K�M+�Q����C!Z�؝���Č�Y?�����h�Uk:����S�`T��G��yl�4^�X�?޻v��7�F���i�����${�K�,�m��,�#t�����s% ���W���C�O���HJ��B���q�����$�~�,g�,a8���-P'��F���Fd�W"��4+�r��/��%���� ����BWh
w#�BJ ���􂣭�͟��:��.�X�#��>-���?�=w���)\�͒x~tڂ1�'&�䖠2��U]bհ���c�+�M�q� N`�:WVRϪ��w����8N��2nd`R�E�,Y;�e^�&%F	5{��'S�J(���S~E�-K�c3w��I�g]*`���"�o֧��kO���5:�$#����	�a�"׏"����ͦ�O�� �Y4(�oPi,�W��.A������-S�k���g,)G 1_x��~3���� `���7��a5�����F��,�	�ˤn-�j�TO�
_�S=�G��$��N�F�A{�h�<��<��<q��F����\(o���ܸ�d��&W��uE���?V(T4 �vJ�=�?�=���@�&���|9��5J8*-2#m4���e���9��r�6���C`@g�OG-t'K��l��E����]0� ��4M�c�W���y�J08�2s#<�3|@���8�>�vF[�0׽[uh�NX�p��_�I�d�U@���W8��x���d�#��Y�S�p��-NQkh|)�U�MJ�J�RR��k `��"�^����㲲8B����JB���BL��m�X��o�B�!�ϑz����1�!M������͗%���Xur���-�:��J��|�]�u�T��b8}��}Z�7��߲��Ĵya��T��_�̘8��ӎLÅ�!�S��*�?���}ǳV�Q���~�P��K:W�b���o������j�ځ[Mq��-ݝ��8��S���+�U{g�Qr��v���r�N��zsw�[��yid�\�.�X��S�L;��'˘LQY���{r� ������,�LJ�	x3�0]R%iX ږ��Y]�%λ�8{̍��)�E��*�����Ч���+�K�m
DZ�-D��䬅w���|ӎ��8�b�0.�,�~1Ȥ.%e�A]��e���
��%�Ai7�g$XU��s+��~�( 9Ѹ�嵔;��� �Jm��j��J�MH��*ч��%^s�F	��8
���Gen�܍�l#I-JHy�Ⱦo'�J�'<���h�����rNj,-��{��A�do��L=��bT�?�Y��FO0��������~͐�<a9����6��oTPǚ�%�V�h0	p�� �
�1ʉ��ƶ�x"o`C�|��Zs�'6W���D~�ެo�NfD��X���_�0�w�ظ��V���{U8i
�ٗ��idn��xG�2{_��,��A�:c�Rx"wo5S�E��k&��.]�����f:,WG���4�A����)�꽣и,ݐ� ���G���(u������������F�����I�!E��{3=T�>���X�9K�b-w��Z��b?L�)�׀�KI��>Hkph�7��DSl��u1��nv�z�����$�;E8��f0㚌	၈VB��z�0	0^�RZ�_>B&���5y8M���Àl���&$F �� ��}1�Dx�&�Y�P~��P�L�#Q�������;�}�4��>�;�~���&Mwe�ܐ�ˏ52��U�D�@�;�u�'F_U��Xq샗Bt�3X;�Yݖ`:� 0��~��	��0�q`�V�����BŚ�3�+�F��H*L[_Pu�}?79�~��lo�xL+�q}�L�P7��A���\����sl���T��jv�����V��C��{���|O��*�y|f�V�������\6�z��j�1q�V����K��x�˚� �frQ��.7|�éoP��Nv�^��o:/	Rp'��w���".�DV��J�5r����/,��(ܢ'� �ۍ�ּ�0�Y�߄y��#uR`#g���G�~W����p�e��Â����J�GM/��A�P��^�l%Y@����i3/L��ݼ7�R����z����<R,}]3��K1xF1\I��Be�~�+͔��j@=+�Ϳ:���g��-��c>�t��~]U]�؄��9���/���vt�_��M���i.D͊d����T��7ܖ����<����
W�����s��As2Y ��vOQ=��m�>�)u�����u���+�mw�:0��sR�����n���V.�A��r&P����4�8Ws��o��3s�Q5�n�@X�:J�ac^������~�@� �j��`Y��'���__4ʠ6�[]���z-%wD��1XI����|}�HҬ �,�=\|Ǽ|����J-���,	��B�����_�@U���3�'"�$�,F�`�)7��1Q����$�����������}�"β�E�V�@�u��-Yф��q�mk $5$�1�H2���}Ԥ�I�$x�pq�2Bt/J�^�j\����S Xj�M��g$�G
U4@�S� �>��%�������g����� ���T[�lD�j��Su��~���P���Pq����9=�uIFqj"��mk��T׌;�1��	ٞ:�f��Z ;����B�a/V#���yZИ�=��\3���3�5�J�)H��^Y)��wLg~�T���(>||G�hʼ!l�H�d��1<����G�����~���X\1h��	�FV��CiF���dD�ђ�D7��(�H�����X����E��CY�ċ�QMi�0��:���	C�|.��ap��vj��t~���Ph�l"�.k�E|��4�k����_�`�� մ�wd�Eg�#r�e���d��<��dֵ�����ǲ@�jP������x���^�QF4��*��k"��~Mh֏j,˴e����
�-��?u.c .r$�Y���_IL3l2��r?����-��
�u`c8¤,� trW�\6�²�]R�\hf4;�"�.�1�����*����s���ІM���\�@��{N?��	�n�~����������������}(M��rj�h���[US[U�H��I�b�(h�mM�WN�	��ɜPC��94}g"}�Q��#v�ߟ�
�����8ߍh�}E1@��(��J�'
W��t(����v��R��<^ûG*���2�n��{�6�g&Nr���A
�D<��?��^xBp#� �Ҝ�a`�����2DTl������������j5��xq�ؼ�̷-�|d#�'�W���pw7�Q��j]8��y�HxR����o��վ�,���QUSN�0l3Q��']�ٴ�S��O����^5�W���t:7�fĨw<i��<4I�d��S�������"�bp)X�S
9a-m�C:�l��r@|�F��㫑�c���i:ib~r���n����3Y��&�Cʓ�-��7P�x�2o��31�U����\-��m`���'���	�:��#u�
��q	ń����$T�ЇN�~7b+���������V�f��CD����(��Nk;�U�KQº �����4�9�&�M��M#���_�i�����Y��qƳ�`*�w~ ��`�aBU
��=Mqk�A��`E���oM�J��GKO�fFj�&wb+Պ	Y
T&�Ƈ�=�D��[)�	7ad/��R�7�����i�m3����쳽P��R#���tC�@v��w�	�^�TX�V�H6�OV>G���͋�@7�5�U��EZOխ{��Y�Hek���0:{�p��&�_^ �鐸���>��$&KjG|X-��@�>h�[�����M x\0S���1X���vV��� �V'�����6�![�h$ ������V��r�/���~`�G�p{{^2��Y�:!Kr}��	��5�7J�e1�q��>����`��|좡8��jp�QQ^^���#��?� �����_��;�ԙ?��.T�2����B�$����\�}������q��FT<w�ɎU>f���%�f�)m�i9��vk3��eti�FE0šLbY��o��*#,�t�`K�����w�E�(�0>����9}W\����� ��P�"C��c\f�'Q�v�������BBWC:�6�>�{��͠�Þ�Wj1�G�q�鮓ݯC+�im� �Q �ZD��:���u~��عA_��$���myg]`l꧑`	F��VAz�����5���M1��9r�F�貃��.Ã9YB�IT
�]�:�?Yk��):=x�[�$k�@�-������0�z�e$U��mz�uFOZ.����L��цH�c�ľ�!����DxB�2��[1��`��>'�[�h�Ǚ�ȗ`���3�~��Z��W��6������̘��H�H����:�8-M�j/H���]��;n3�!�q?�>�Z͋���������MP/P�p�񬿧J8���G��X�q�����@�Ӌ���g{�Ȁ�.4}�X�5'#�{'�c�F����t=Ʈ�Vŕ��9�<h�?���IZ4S�ƀ�]�g��m9�&���9d|��R�+�Q�������WG1�41s�[o���j�*z��WD��
Ǹ!�	�<�������Г10@��Ƣ ��8��Zl���X�O#�V2����ψ�)f�h�2X����q,��ѱ���B����hWR�i�9��]������3��ױ$9(Չ)Zl�E���p���p���0a��&��S��o��!&���H��#=�6d�ypc-;F�W����I�I|+E�K��I�m-J|0|rW8��7'*S�>i�J9?��/o��B5�U�z����1��+tq��|M�T}{��b�"�*|^8�:���c�����O�JE�U܀�0�t}.�K�#�,��Ä��v�z���e�-^'z[��b+���N3�X��l�>;�EKK�GV�'�|Vq����(��َW��:�P��v$��,ҫ��mz�|�:U�4ZY6d��̫�d��G���2F&x폧����"��{������=l���vVoWO�Di�ÿU.�g�/�Jaȴ9s�4�!� ��y���A�zYy�0RRl��X�p9�|_h�J��E�&�ǧ��eRu��EK�TT�t<�=��(:j�Dq'N�#`�< ����4�n�j�R��E'Y��^�
:�y��{�����$&'p�+��O��X:���H�a�\3�;x�w�,|1��\��Hr��qA��������v��*��e�$j4ï���}���b�>����^n�"�����F�<t=����шQ��������.���=]���`��=�PP��W��(Ğ�]r���en��Q l���̵�����3G����w��Rq9�K�����}�UAxg?���a?�U!��k��<�A�S�?*� /-�:k�G�� 8&"&K���۾�˞;���"�/;��m�!��?tT2��y���*��`I��߅6@C�v��X�ڭ]�Ş�|�,��L�Ҿ����m]'ŝ�B�ͧ)����5~�|��{�1�{��!���u��ʽ�jr�U[�����l�,rE�v���r��gѨ���	�vkcW���~T�fz�hN-�m�7�Q)*0q�w'�`Q(���\3@�J�-[�僽lNM��4b�ߍ�#W��vf �1��q����G��uO\V ��5u�����6v�ǰ�W��l���W�t@��24m���-cS+qh��kܾ��ŋ�����	L�^�~B�.�b �5)�帑�>�>,���MK��C��|#��,V�A@%~Q/�3�׃A�\A-Y�?Z��R�,f�{��@��0>Y*�w�CŅ���1�T���U��������F0Ta��q��ʍ�o�����	�9R<���6��?��܄Gh4���0p+��������o?Y�A�T!�\�S�z�;ÕW*<�1l�����������Y��GS���~�<o�Q�0�R�f`/I~#����_�A�9�S=ROޯ��}s'ǱZ�ة��9Q�=�]i����O�E~��QK�i�W�-]��D�9Q���Ev��K .C�J����Z5�
C�%��x�(�����@����+g������ֿ�C�bB�z�+�a͟��18Ioa�a�{b�OJ��/_��)�p��x���q_���)�D���H�*�Fģ(��n��:��=H���u� �;�T����Mk�^&n��������	]���ع)�e���[�_;G��1W� +5�Q3}ڗ�r����XK��c�?DT���i���7nUoi�I�R�2���q�%	J�J�|��Tߐ�C�it�>V��dB�8�έ��y������S�L �.o2&^�(OG�v�(��eM��~�87ݿ�������5�i��2��n�g͑ ���;�ҁP��e��R��x����`�P�0�6Lt�-�Lt$�M���*,���ݦ�.�f9��\cƥ�{}]�ߜ�w:�u���Uڙ�R�8YY��M��v&:n�]���M�&��4��?p�Q��D�?��x�>�#}}Xo�mAN�1�#X��/j2�F�,�ʃO\��t��TJUe�u	���q���Pj��UOG�%�&�#?�*�]J�cWM/;e��.@�Á�gM����Y�N`95��	Wy�ܔ�:��	Y��&u�1y߃{J�'�2�O;4c��U�Ų�)p��B��驅���#��-�E��L3�M�{nñxQzz��˕��_����[`R`�� &U=1��S{�R�fc�9b_Ioo3�H�\�־��u�o��8��Jk&�;��L�-{R���<�[%;���?��9<���zc�q6j��6��m�vۘ��ƶm�jؠy7�������d��[�>g��Y��D���&R^��W� �B?R+l�Ð�w�u�a��Uֆ�X��f1���j�T� l�l���	��ʉ��4i��c�E��l+�)@�]V��r�.�.��3������:ibDtm*2ڷW�:�}��Q���lQe��Wy���˽��x�ώ���_4Q�(n�3���:���]�	W�|m_8v����"�I�>�;N�e� �V=��O}�=3X!���F�P�@MO;�@?�l���:�5y�Q%�ڏW���Oi�S�ZO��ɦ��R�ߨB y���j_+8�*�juLrj�5[�zԆ�퉵S0mޤ�Tj�C�vQ�\��������;�FŌlv��W��+%��t��_�������������W4�t8�-�L��P�!� X@�r {�2ב���v������yĘ����o���!]Z��~vD���F,��FN÷�$|��-�>$RZ�~��H�w�4fb��OD6'�Z�Zj?��@`�jk|��������8��f�{zNd�2�������E��{�ȁ_���Zč����~ =��/;uz��1�Ķ�9=V�I9���29Q�)7�J���7��2������ܨ�/��,�'�-��$k5 )4���?[h�=sk�yK��S��B?-��+R��wi��%��;��x���.��\�7,��Z*'ޟ�*o��,�1�2x� �W�4�:Hws_K�$��;����L��	��yK��v�S���չ���I��HZ�(�i��Ռ���W¾�_h/�#x���D��T�}�ǽs����苼~�>j���P�)���A�v��r���y�Jj�&5v<�0[ۍ����p�_����W�-m��9t���5>ˣ�"��X�;B������wE��w}ǽ�mŶv�8�4���f�6h�-��T����Z'�qJ7�,�s%3�S-@�wP��~~]�^�&e}�2<8X�;��	{AP	����/��=����Z�j�f����Oz�M���~s$@�~KA�Eψ�ɯ��`7��7�Y ��N�j����� 3���T����ᖻ�"|�x�DR�
�hr>��tG�DI�8d���	!u���+��Ȱ�8�U½)8A,}�W�Y����;h��5���aP�� ������+pYS���c��
���Mg]?��o<�����-�3���������T�V��k�+e��Ӎ�J���_�������ޔ�@)6�'ً����j��� 	�ɫ ����CN	��+�R$�.��7�{��������}F�׺����7�����u�����C�fZ��3*��Ʒ��*wO�Dw��v��
��� �8���i���J���]�{~ m��y�,���� �`2�O3`c�
�vsO���&�b^�=VmG��'��QǹߢQnS[Z��,��!M	��n;i��C�k��i_m�myG� J%K���w;��K7X��3я"���Z|�_(�x�M����3����uZ�v]�%��@�J�T"����,�!�,+����K���u/-*���t*��a%ޟ�J�[�v*r�G:/]bk��i���O�6zLiM�V�����t�4�mG!���Ԕ������_3-T'==;�Ϡ��%"��R��Ǹ��V�P��!��>�u�FS��bi�������}�k�y����u�z��yv�y�F��+j5tn[�2��Ea�n�,������3<N:Z�O8�\��z��_��KL��9/C8�/OCt�|H���t�)0k�e��r
\��_��?Ԗ؟���*�,�A�nz���y��� £�ص8��{Z\�����-�(���ӿ����d�Z���7����j��f,^`ÇL�u�2g!"����n��� v�^g�)cN�R3�V��C�/G��>!�A��A�z��+��1���ȿ��,a��CEC�^po����3�~��c�+�[�.�������͐H�u�ߘ~��X�#�
��Q�� ꭭����%D廧�r�7mSg����J�����A�t4���˂����^��Q�J����ӓ����;���fBٛ~��I֛��"�E=6X��~������m���;�Nk:�bt�[!{눛�T�R�����`9�h���,B�̻��|ғ]��;�/+���=R�cI�x�o� ����a+f%t@�;U���/�S�WTo�L����(����ٹ���N���[9˯�}������R!�?ɩ7�����-��{/�z\�/K�|��X��}	��eT���{搑�P������E�9u��]w�r7,C�Eqn�PLj���Gh�����x���Q��BxUVZ?�3���_\�ϭ!rT��'!���ż�������rY��у+��7��iyx�T3#�ӗ�o	��󰍜،�H��J�p2�W�/���P�x���ޏ(/M ��O��R���z9�� u�~���u�>������AK-p)n��-����t����6��sj������.:���*<�r�B���@V3�����4<���㺪����ʒ��m�H����O�	��u�� j?�J�|Y����`�l{{,��	<�U�!�&���RWKI�;���<�6����x�ʹ̎�ڂRK~f���;��s�a-d�y|3ל1�S���{�^�z0WΔm|\h�г��p���!��Wpat�P�ӭ�����~�][$������Hf�]�θ�M�-�}�Cw�J��e�;Uk��j�e(�
#�����Fm̧@c����=|�5ՙ�X��n�^���Zs:�W������jk3��ݷNp���~�f�<��5%X����a3�6�-�O������_��������I�f'-�a�r�j��a�B�x(Ե�5�~�'�Na��aG�6L<�M�N�O�{b�`VY���@�郟�V|���/�pѥ(�P6ђ����9������`R	T��/��स#��q�Z�B���9����ONp�^�O؈f����@�j�3{��HE-iL"!S�̫l�bס}�V6��3�ڮ��Sm:�VK�0�a.������<nI���M�Ӓ�f����sz.�����'U�y=�$-�� T:�.|0:qwbMN���Î�4��������y�g/X��������)����S> �@�.*p1�Z��C�%}�\I���Ѽ���;u{|e�U�ǶyÞ&u���)����F�m�IQ`�J1G� ����-�=?pK1���❮
K,)Ӂ�Vף	���������VR>�Z��n���mK�C:�g���}*ըz��9�@��̏Ef0��1_��1�j�.V���{�U�Ǫ{'�~V�nt��]���-� 5��ݒcm:s������~V�}3���f�؍�<y����Dy4�B9T|��Ҽ����69qOu:}�c*������G#P�9dRv�z�W�
jLY�$�6�RRR�?-_<�8���<��Ԍ��M)��o�K��l�N0�GtW��[`ќ�7�<*�"Bt�}�_��=��I;h�����Zlnd�@��	��r+*�د5���V_V7,a�>�^u0 ~Ճ�;^���e�]�q���������gϦW`��^�'�J!�Q��Q��UBV���&еD�r�P�����<'=~����cS�n�E�]h����C����B̊I^�P��[n��x�p\�b_�
��kcz|q���`O���X��e��E���E�iRw�U�}
7�5��Eu�é�n���0d�^�g�{G���-4�;!%̈́؞,2V�J���N&iPv�'�扥 �HD'��J�������){��W<��^��f�L����@�m?�1^�9:�~�����I6�;�\ai3o;//�k�,4�	���_֮��q�5���!66H�)�e��}۹�&N�^ڐ��_�u-���"�� #k����tß����,��醡�l�{O��}-�W�\��%�H���qk��À��Ο:���fB�ą����� �v�=3M軎/]/j�G��95r���t?%��{`�/c��&i����Ssc[,�(�k�%��؄�����MD 	���LL�9����q��]���������m3t�_.�[�j.�,B�X�Ł�����N�s��׼�y�)ׂ���E��Q�V�Թ_�=���&�r�fZb��Q:Z�� s��e;� �Ju���RPz�<��=r�ֆ���s�w?����-8�����Z�M�?e�����RdU��-�~ߣ�gs	(��t!��=g!�V��%SY�G3,=|�6X�>{��dSn�D��WNO��8�|g���qO�j��
UK
K\���V��G�q#�F_ �ߞЫ�4�
���{�*]�(�'�Rz�gqW���w��o��-�̉
�$�op��jp�%l�E*ްx�Er�\�=�J��"�����3��=B�F:�ʠ��粺��b��B'Zo��6�Q��{��.��%�	<mLZ��)w�@�_j~�P��W�l�Ѓ:Zq�+���.X�=�)��\�4O�ŋ�C�w/�4��,�y��j�7�M��.��>�x(y�e���o�	y�֛	GL:bt�s-����eM�Ġ�.�*p
�&g�	�h󳙶�{�ܠU�N�����7o��݇�����jOW�1��J�Kx/�����o�Ÿ"T$���Q`�C�`�̘���-j�%�`z��P�y�$�� t3��]ʜa����}�RT�E��2#C�Z���Z���˪s�ථN�:�(�~�,.s^or��o���_A$�z���+�S�N�����|�6Ƹ�� �]�zx/`�
�~����1iU5=�+����\��vbzS�_��a��f��ʠu%�8��ӏ~L��y[����9��z����I����)_��v�:������}�a��!�b��P�Gk�ބ$��ţ����%����
��f����b��w=NVa�2��Ȼ�9��v�ѵ ��ng%�r*��ղf��2k��/Dܷ̬���F��|&�ِa�B�n�}���\��8ƪ}����m3J�K�,�
T�<���Rv�K�e]&hS�_&Y��ś^r4+�{�B���?zХ���7ƅ�Z�B�P�n�f3/�1��b?>���P;h�2QY^�]�4rϱh��7�)�S3�v��<Bew���sm���S4�|�f�Vv	�^Z�ؽ�}�����5�~�_yݺ��la��)�D?�WD���9��l:��Mp����B�%���yA0ى��~�`��дV��A��a?9�C����8�I��҇섩��O�'ߺ\�|A�h	�g�ig�O'n��\��k��U�-�{O����Ll._ֈ$� �����n`�\c��^�`�_	��;K�Z�%�*4�B��+�FH��'�z9Ga7�T�e�J` �:9[��*�^��%<5�S��(���3k>$1{Rl$<˻�[�m���<�{�E��sdU쎱:�T�&5ڭ��c�s���9��;�p'��	�~O����#V�+���h��@qm��K�����8�̻�3�`B�{��%UG!�F�Ėee����^�~ס����N,�H����͒���/�,eLx�%�[蓼謚f��D�^�ƿ)�G��i�dϙ����E�y@��ʅ;XI�V�wj)�jc��ⷊ�����d����s�tuuݡ.my3�b�D��Nm�Z8�Y����}5+��x�;6q��q�|L���(�+Wg����+�/q��p��d�}�鐥�a��p��Q���WT�����*}~�i$f����)�J�8X�DҦ��mu�[�{1x5�$�y'6���{y��V������&�H��I��u[�=r+_����wfn�4��4�&��v��S��H|"��bf�l�b��9c���-��0�����÷T#�>�[�ʯv�6��亁�Hω�S1߽w���]}b����B��8�X&M�JG;2��5���c��������q��h�g�I����>6�j�fէ&\ �A>g%�O�R��>p�ǸV�HY�`����̶'̣��;��0p�#;׊�B���{;�X��f�E:�ٽ_v��ǩ�̃�M��_�yR̀1v��x>ܶ%�J�I �G��I��ۙR���N��.�"؏��h��ef��>Q���$�l.o�\`�3ٟE�|+K�nY@~ǚ��}��=;�����>�$�8H��.����~	'��ej���Xj>��~����x��{�\��;@�^�k���=�7��T����.�p��3M���N|�AR��LT\�54�
s�]�C��e���(+��%4�F���m��:|�(���Ѻ��;����n�����ϒ��4��|%�)������ϼ>�:.�h�㺲�ZͰs��3�j��������{��b��P�Зb�u�Ibo\F��(Ip���󺺄jv,*z"H᯽:�x�&��W���mB�EU�;����ݛ�"�SǦ�7K^��Cm��zw���Nx��Q��03lp��$��G[�1zn^VH�=���[F)�n�`q����qG�9������w_������c�n�v%��N4��Þ���w�3*9[�Gj�G�_���i����ι=�Q��5#��`ăe�}_q���� 7f�/�w<������k�r���>cC3�t�9���9�o��u���bϢ�1V]ahl�3�i3s9��N~�����){=�(⡮���#�~��*�a��F����M�G���Xt�Ø3�|�ǌzG�r�9X�͑��CN�܌�~�R	#�	R�xT�'@j�	������V��Չ���%�H���{ͥDB��8ߔ�1O���_~UZa�&��z���x�x
N��H��%���ܑ'���D(u{�b5�LV�a�����s��B٘E_�*]p.c�Ŗ�y��כr� %���]�<l�o]%�'��6`s����Z��#=��2A��>�e����L���B��@A5Ab?.Ϯ�2ĺ�b�P[�xs+'��R����MoIi�E�ͭ�C�/�'��@��		
��转��{z�P�o��,&l�;��W�s��0��-�3+II�A�L�H�����p+����"Y��]�����˙�q�T��h�.�>�{��F��������"�kk$�L[���$����>(�h4���gI�{ĝ�ȭrjh���ԡ�\
  �d%fbq�*���0VF}g�� q��J��n��I5X�o�&o�QC�A�0e����:����-pv�X4�uN�/l��� !�׃[�V��4G�R�g��r|��܅u���2�����Ȣc~�+`�牀P��_̉���WӞO��%���xe%ά{bV�X"F��&��%�wS�s��Ɔ����{�����pb��!��W�]'��}1�%Ѓ'�&aDBE�'��_�B�d�58�=��W|�M�G���0������x6���FHO����I�pUf�j�6�r��l,�Zq.���o	�X�y}��4��Xe5
i(A�A.f���$�Wbزm�[�J�ʤB��K��=��xȃ��w��;%!8]��qT������❯f��.�g}\��7�b��)w�4�^�}ї�>lh�
��R	V&�T �w�'gm&�4��Er�]�����ڻ��r�dh�f��D��a�y��uJ(<��z�Ո맶ȋM%#F�����xĨ܊��i����t��UB�� A����9�#���9���l	>��{h�����>��r�a���v���	g��� gg�{�/NS!oǇ�*��qY�$,݇,Hg!��U6)�kJD�na
%!W��C\wH>��ca�?��Nǂ���kz��� Ph9F��S^������c2�<y���(�-zm��q�6+O��Z�y{
]��G�j
�jD��'�ά�5~-�J'2�%2;�SQL��y*�.#��p��)qH��� ��bK�B޼g�\k�a@i .b�,�0�Nt�(�s��Dj� b(L��T�ʖ��y50����t��}#"��]�������1Vi?���4���D|rn�-��X�]FԊpE�x'ki3ڀ�fh�C�����(�W�埣��x۳�w�Ӄ:_��bC��sÁ����oRY��	)�4N�t��X-r�>ن���fP4[����E�Q����H}�7�&Xު�)��!�:k��,��KC�,�Hu	/����򀀌&� ��a�M��SY|m��y�ƮT����w�� �}J^�R�����Y����1�fΔI��K����M��œ}��d�.����ӫ��@,��Q֗�_C���b��w�a�o#siJ�i͂���S��'6h�ⱳ g7)���p�&/ ���`s
��<܎0w��c�p0h�h�5Qi_/̸�.N�v>��l��M�Y�1	�Q��u�/U�*���� �7ak�!x��E�wB\Ȅ���$TB�-?�8c�z=����ZD���B���A�+
~�Ϋ���`���
)�3'p�:�k����N��bݗ��u��}����KN:'Q� [��I��k۴�
�u������E|)Z��y+������"���W�q���6jl�7��=s�^H�ڠ#�r�T����B�{���:���H�z6tn���ED<dB�X����}ܹ���y���ku�bSP��.rE��_Z^5�G�x�̰��W	2����6i^!	�)[�(/�Ѹ���� t�t7�'�>��zIX��y5�[�uW��"��Wn��屁cw�C7�Q�7�%�~�������������� nA��g'�0�1�h�mS��3۷���.�A�N2l�՚�Fl��@f͎�W����8�u׺��q�f@��%�:���x\���d*}�o"�������SL���u��:9�­��:NL*C���ڮ;/������������[����B^����a�5�R	�.?���o|��^��b�$���h�m`a�*��H����PpX���ۦ�g���/�m���b<h(���B(�؆2x�輹^s<��u�'���ow)Tc2���;� ���I�y����K$��yEz��(�qY�5�11�oH�:�M��j�B��7�:�^��k+�g#ˇ)��,�b�Ȋ]��v�,~T�3��<��~��r�w���F\;��﫟�ܝ�1���!̫�S�J '���N��NO@��mZ�q��%r<�Oq(�&���fki<qdV�3�$C�V���5Ig���Y���Zu[�	ў���®rZ�wm���^�xe�����U�Ó�7��ԁn�)k�ѱ^؊y�vm�^1��)V\X��Es����)x�
RNcu7*��u����ő�'43I��b�ם2�}F��2W�y��@<�ic����>N��f�2Y]��Cz>B9��jP���bW�8��- H�D�
V��VS��G�[���~��s�/�����&�^��[�鈘���2��=�� Y_q��DY�Y���G6��Y���QM��9�(����'��9�xf/U� u�.�Rdk��m��k�R��,D&(���]�� H�[��s�
���O�__ �o����
�jxQ.��n�\��]z�s�@5�]t��ۉ����=�B�{���g5+:�<+�[�g�Z/���o�t�T��O�	S��Sǆ������j~K��G�W&[�.��q��#�^�ǩ|��OA�5�� �[G7�&�t�#�yW���Q"�/��{�0�龖���JS|d@F����4a%��|������zzA|q*D5wat{}~��?OωjA���-2h��6�� #�ɖ�׿��s�H��_�ϗ�g�B���/H�F�>'�I���$�i�@���7f�@��jED�~���"��1�qLX� ��R����~��<�7Wb�+� ٬u*��FLC)�?����r�� ���	E��x9��>�;f���a�\m?�$�a)����V�|�Ġ�C�/!��pC����X�B ��E�"��JQ>F��f3 ��cu�p%+~�2|p7`�J�ߜ��~a~�l��;�R�ul���6���	�{�D��[���|��-�Ue�rBAB�A����0خ�K1s��4$ ����@{�?= ��NŃ��~�'߃`���qa#X/tTJ��1aP*�JA�+b�m� B�	Tʪ��>O�[��_��S�<�b�Z������c�m��::���B�}`�ً�.1Pc�V��jd�b���$��|E� 1ټ]��J4ɺ�<4]�ܺ�	@
���@d�7�t�v�����^?O��tR�����ܔ��t����� 9Sxk*[h�����@6�ȣ%k�F���t���O����f�C#H��kSx6�����ܦ\�D�O�Ɲ�a��[�K^�D ��1$8��N��9�GZ�O��)��X�Y<b�V�ύz5�:�gb.j4�h�`�����`�d��"e�ɣX�7?�Y�D$A�CC�viN�2�n{B8�l����f��4���E*	h=���qQ�Z.�� �!'�w�/���F����~�Np���m�������"��w�_����╳*��*v�|=o_�=F#����0�a
8�4����i�K�é�1e^�4`�KxLj�so��K��J�ߖ��.���JǨ`�

��^fA�������7���-`�$� k�/�'�)�P� �bG��,��v-K��ϵ=ۄ(
o`�1q�GH�]����Gݔ�7�i˛\��
�
���GvE�s!jB����֤�v��ω�&�CL1�QH�F�_,d��e�΢�B���L�Kn�~ɐ��n�%��ZO	�9�)��]�S��r�J�n,E�J�@!�EI��	�h��K&�ԈY[^j7�ݛ��!��,s�4Qt3M�U*��:	�>dt��_��&����$-����셼2ߙK6i��6qk�h����\��_2n�Z3�<��+����'�Gh�����q���m�5)ȸv%y��$�Y�/-*�>��r;���N�K��zc�:�@Ǌg��&��ّ?ު�����7�f�*�fjܳ����y�璡�􏑙)!��h��l�AD2���k�w�&����1�/�P��aCd�� �@���<aG��	��?�9��B��>�ܢ�Ã[��a�9(�,���:P��9@��	��p�|�z͊76�҈$PD��>�B\�2:�w�ȵ��K���G�۞�!���_i5wRYԣ�m ŭ����o�B_l�5]�Ԑ� �&��m��3=�!VZ�cE�����ѓ�b�B�Y���${]#�w���"�e����F
K���JVPƺݴ2�an�J���1|ac
��0Y�H�H�����d�qx[%T5G�� sX[��[�*�(�hi��k[�;D�as��m�
M�j����?'��a"(�@�mTҘQ<�.��<;f4�g'?B������	'X	��!��Q� �4&�)(�O����٘c���!��*eJ�%��dkt#Y4}6�H+-qҺ��f��Ǟ~K4Uq0:���=�GrZ&C\Ȯ���K����u8	Zˮ���m�I�IU0$�N�^>\��aYrd��"6F���[�����9����ԛD{˟н�KcX���~�D��78{;�3�Q�&3_��0�w��cS�Q�Ĩ$^H�!�s0��%<�K����
�j.5���c�'����+��~����g�W*��o��,Eyq�@B����/�_I�Ӫ�i�g��c�����?l#ϐ&͈��뜕5fN���M�\�t;��z�E�ZrQ$�� *�؁�e��(�#�l�,Y��z��=^��4y�����3д�%�ޏE���8�"�I%6��}VQ�9�'_xh�� yD�Լ��O������d%<�:��Ơ�~��ď""u��X���*������>�DYW�GN�$
f����	�ec���;.v'��㺽����D��Р�A/t�W��&�M�#@�"R4FN����2�0�ra�p�j���Ѳ�I��0ʺ> k�;[ք��+0r�FT%(�v�-���;�q�AQ�� �!+�8*�"�6yj��:1&�K�,Bpq���J�FBM�o���δo���@p�1��i���<���DSB|L��8LR"�ABw��~]�J�vh��r�,�խ'���G�QQ��Y�%P�
����k��1��Z��"Q	�Nz>�.q���3FJ
ja2���B�(ѣ�=�$��s�0`di��pm���2��+����Y����2s�J˓vmH����U�aRR0L�Ӑ�Z;<}*�����^�ƍ�1�Uо��J�c�2H����F�Qc�|��} *~�P	%��Kt"5�+��I?�(�SP�0|�]q�>2j���&�|�!.w�� T
��B׷ �Ȅ	�S����"1�9����,3��{��>��	� �S��Mi�1�� L���7��5)P[M���9Gy�a{�B��¬Jh��Sy~�8+�͉-����>�@�!a�7#��[�0w�(��O%+�h<�)ƹ��ɠ2�mO�����v�(#��ݘ�?0m�+��|2c�dpt�y)�&�!H,�s �7@�hbz�¤��t�BF/Ch��F��po�����K�.o͎��I�_��p�BE4Nq���q������A9m?���H3����l��?%r��o�*J+N�*J�{�O�8��R�Z6�"	��͢�$G����d���+�kg�
\�
L�n���Fx`xt��+��ݯ�~��u�N>�.3hm�)�CY�M>O�]^�> ��r�)@�;,͗X�2ǡ*�Ƴ˸����rf
�&襳ן�����%+�˞�:k� �4�y����Z;�b�Ve�����sT���Ul��D�<E֑��M��1�_[[{\.��Y�'v�$
a,h�5#��5!�{q�dn�{c:�]V���i�|3�(AE�R9X6��ƀ��"Θ��6 -W�D�����%Խ�ݭ
�W��ȡD�"���KA����[�K����U#�/Ն��+��^��re���#d���ö�m��2����4�_6��_���
��Yp�{���	<��������Q�p3��������qF���9� ��k�:���y%�J��#`�:( l�'p��R��P���<��^�M��UK-t8d��C�����_DO�6�5-2!k�����p��0)5R�y�M|�hCu/Z��R��0*Gv���H�ly	C�3z�b��A	o�<�a� G�:�u�b��]��P`^��񋅚��%5G�9��?,� ��tD���mb|QvN�&J�p���:�5��I]Y:`�8�;�O��w_.�p/o�h;�:x�*s�U�^G�l�p���I<dd�?+���Z�x�mG}���;\۹����v�X>�׾/�k����@0��6F�m��g�/��u�mϼ����Ȳٲd�{�R��;�Y�@�M�$[�~� )
�<:,�d�d�<����^̀T�$�"��{�,D�,<�ijv���(cRm��3Ε5�H�fƔ�L��O8'����Z���S��rc�E�ͷ]��H5ܴj����F�mMހ+�Q���23�5�������'ohʆ�RP�6(�E	gB��B���M�s 4qH�T�`�D0`L�>	�
��IG B~���Qc�!@�v7 �
����!vb���_X��:M��w�����Z�4c��/QM�Wj =��ư�jA9U_f�@9Cy���I+���P`����|hc>(I$��Yoo�΀�l�x���I4� �싸a'~ȝ��'C$)<�Vѓ��%3W)^�i��b:�O��_i6���)���}p�Ņ|R���
oX��-���ޚgH��� ��pE�J��D�Y�@p�ƕ)�Q�XENl�h����rH�`k�5bR��9-E� Ր C2�8������/X�C��]L�
�PqF餝���k9ׁ{{��>Xα?{�׼��N��$>��� �Uz�+㯞b��Z���#+��]c�ˆ[�2��y��?;]����=4��ǯ���lIcS���?u�y���{��)x��S9F��ո�	���,9�^���`M�
 4_G�DLݴb�Ǌ�>�B�ۄ-GfyۇZQX�!J�B�Br��~�$�TF'�e��<\�p�T�7�<��%�y����0��J�tz�$��
�+?S/*x�f��ş�%�b�8CZz��;\:/7�Ql���]�X��l<��0��;q1��@X���f��Ƅy���X�f��1�'k���yXBm�6Qi+����#�Z�
���T������\Ï�~�8�*Ĉ�<���K�s���.̟vI��l���2=D���
Ka���V/�4�*/C�SgoT����7Q�C�]�;�ø��l�o�~*Xf�	�G�/���=�:��7��R�o��a�Q:��mc�x��f�'֪ż�����3H��Cu0��l�J��~9��A0�M���t�$z3�gG�P�(�� �ܻ�^��`:G���nژ7+k4���L��	�b{KT�j�F�� ,������ߥ	˫u%��Cy����:��Ǎ��'�c���c9eS.���	�?D����@�8X)(��R�,Ov��N���f�<0��
e�������F"�z{��Yp�>�F�H�������:b��5^�u�S����1.��!ڢ��G!a�9�B���N��A���j��&s��p�kM��X%x2K�ӯb*��W]P�c���d�� 3+��ε���u��8`��ວx[����b`�!DHQ�,=(����j+�6��������/o4���btF[�6�dm��
?9B >i#��;����|�psם�<~��Y�t��C�A�=B�o��/	j^�I��j�yN@�
zr�$U]���{�a���Rm���h�6���^�wϥ#�]�ؾ���@{=�=:$AA�q�'���(s��W�u�%8ǽD�1{��_�fl��9I��҈"�M�����jъ��6�p���{ n�[��h1"�z��$���67q�AU2\=m��(��,\q�����r�e���ܸ`]�-i+	�9u5$p�^'��9Ӣ�������ӡm��F�6t����v-���o�_�惇�����\�u@������m�D����W[�"�yد���{B��$�������mO%��l7�VW����BG"E�ΨCv{�h`Q���4_��wx����w����]�0�Ed�����M�oS[�%.j,�\.V=�8tz޷��k���*/����m3 8!��a` �xrN%n>�������R2�d"=�L}:ZGV� ��I�+����|�1S���O� �O��5N�|���r+tnFM�U}�:oPR�3Ћi���R���z!^������NWomh�����"D��(ԌKx����Gg�'đ����t�dH�F ��=�������״uk���J}��u6��Gb	ĕ�5���!�j�c���}��䶽[���fΞܭ��S���wG7O�(Θ�^4��m���	W	�ɭB��Cf�	�F���*j��";��ѻ
�������+y���sHF�kśH��xF(�Xh7b�^V?���-c��<Ʋ�9n�9��I��@���YO�1v/<��hQw����)��А�}���;|4>ɜA�������!'C-�9ݺh�7�O��j[�R�Mer�r{T���Φ@�M��Pi� A"'j��֝�f��F��k��I�;0HH-���%���O��*�04G����Ī:C���,E�34����y�.�0���ݦj�N����e8�3ނ��_i�UZ��V����7����A����2+p$)�H��v�S�����{�̸�[�U^w���^��yN�"e�m�áM�밦T�	� ������J��������pf�p|:�W9>�-�6��4n`�L �ޭ�$����'�1�L�)�8�un0Xނ�2Icⅱ���xLA���YA�zش���`�Ҹ-���߲���u�CV��SYcJ�����/h[�v|�n�4�1i2J��*��"/]�y�'<�qQb���ٵ�ZT�@M��G���&�}΍<7�sW���5M����']��{�>�U�E����n[�^j-��t��o�v�ww蔕X�\��_h�]�L�vⲾ�t�;�~,C|��b��=�qb��h̾�2&%�HD��9Lgc7A��Ch2�f�c?ݪ����dԸ�}�Fʄ��*A}��wIO�c��-Ěf�8�o�3I)��ʎ�(]��?o�5��+�~K[�Cx ���!n�h#^=Gu�����>s�n��I晃7`�!�]�$�{� Q��{���s�����t]=��A�P��?wZ�v:p��^نn,�����'���=����f��e��_/���#�F����^�C{!��6�6�۸%�^<n�l��aTv8��F!����}x�hva,��ЦZv�0�����ZK�*V���{&q��=k�b�?z<�����Yo��E�.��n�5��C �wwwwwwww��	�Npw�[~���{U�j�jwg����{�=�g��?�M��(0yK�1�Lv��*u��E6h��MuT�7�*Ȯ�|ȕ�Dl\�G���.w2���-S�q� ~Z����|Lgs��n�ŷ�:k/��G�{�6�	m݃�Kqs��K��I����$�O�l!�B#-��ă�j�y�bP_�a��.��K,��d/l�2��6�9�Qa�㉜��U���/h����l@�%�=*ZK��1W��V�ċ��2�����xE|5��<���)�-�\���=1��}���M�9���k�c���E)�7�V�U����N�9��Ӻ�_�l}H14�5�7�MU�=�8m� -�T�\�J�R�-tA�^�\-��%��..�/i$k�7[-��<�Q�
=�2G�8�����+�>�?�{|��(_l��xU�辆LR���W�����T���@�׏�X��0^��lg.x�����o[jp%uH��!��x$�S��1z�p>��ce�ٌ�k�`�B[r�8��Ka�6kFuD�����.��
e�*E˟TK�#l�D�[����R��Ƒr.� ��Qbv��*Q��P~@��>�d#��yj�~a!7���&�wܵ"�q�m�ڮ:Hg������N���m��'l��V���G#��%dR�呈�㠟�b8��`�̠�Z������Έ�9q�ݎeJX�Q�&�u����au�#t �>�P�ݫ�G�����ި�Hu�N��܄�]<�X�ӄ#�d�ڋ�����o�yL1�S�@Q`r=�3;,rH8!�� 8�,�ُ5�٬��}S���4�,u��^�]A%��<�x�캺N��x_���V����~S3�=X4�`�j{����'sm����m_1��H�UB��Բ]v)Q"��6���3rLr_��p[��p��������BK!�&�K�����wخ�Ko�ٜ���FW��(���"�b�s5�-֢�S��pc����r�r.���ɯzX�2���#��j��d���M#���"H�#��U�Fh�H�ZkJ�_��ߐ��c?�Q�;M��=�y����>"D>�y�� Q:J&�F�y`o uf�L������~>�~��Q 0����͎�_�+����bP�C6JI����T�q���n����u��q�m��j/�?��l5��	��H���a�z�)�q�Rf���iR/j1b�#��/�ׯ����C!��f}��4'��亵;���^d�/��%�X),8,����Z{f��IL���)�����Y���.r��[o�����>'1'&�0y�>���ꕍS<,���?�B�VyJXIe����U�`%69K���t���b�PluUsD�����	1!:���I��� ����_s�;m�3q���X��,"T_�.->`��^�v'���.��Vq������y@��y�0B�e%�A���X45&����iV~�g^R��WZ���t8),��$Ðӷ0ҽo~D�6"�����O�-q7LƓl�;��?f�c�ٝ�[]��[U%�W%y��U�� ��<{�V�ǣ�/J�!���.���|#����kp�rON�}��"3U�#�Ms���|�G�r%��\���	���Y����^P�G�%���y�|Ք/v_:��im���{�iV4].vZ˒_���yc�
�D�Zz3e�`�vY"�bʣ��9JB�E�<�H^�F��k����F��)�@E��]jf��(�+��58�'��'g�R��������Wヂ��?Fz.X-C���N�O�f�h�X��H��DS�y>��hbv?��8��2���g�i�o���)ے{�B5���ds�8 ���)�8b�\�U��|��a�J��7#\�I���C�1.@ߗi�M�뾬A�Y�׉�$�d˟�zܪ�Hߦ
EJ�rIa��J���b䎦�J��a �F��Z�ʪ�-�)d��5�(�W��JQ�P�͆���uC"���G!���{��E�f ��� v���X����і��8vU�m�u�Ʉ�󴡜�)���ΰ�Fm{BC��ܿ�e�?��%bSa���;��;r�ГqU8�� �2Վq$i%��qj0�<�@-5!��}��!�H��U,ۛ#�A�/ʛ�n1=.*����]��.�R�ٕ��H�v�@��b���#��� �����'v �%PCLk":O.�_�7!M�p
�(�h�s*��eH����p��Xi���D� �(�h��E������[R��=c���%�oPzb���b�9�K��L�d�-=�^����b��@E���T�ͨ������K������24�M��
-ǝ�,����o�B�.y�Kvv��8F!I���;�1���{��q�.�+��z��oBZg~���*\�ď��V�76�X3���#�צ�[���Y)+��"�Y�(̎����_�Q�u.��Q�b�:59�jM:f���#����0�����J_*
�xK� �$�`Ie�Qq����yV���f�"�#�0�b�#X���_���n���y�k�O��	�v]�V-��j�S�rf3`��R�ԚY �耱��BN\FR�D@ӎV��]V������ËVR�+�Wa#�Z�W�����v�
�g�3�Mi��%e�'� ��Pm��M���ۥ��������F�I_pI��~�evX�4x���I�ƾ��oK<�F8��Ҵ���������~�feb�
�0�s�I�Q"�}�x����e��T�'�wZ���~,����u��l}oh�>v��������2�bñ�G��{�acMu����ULw*z%l��bsd��� s4��7���ƥ�q�ُ�&�[{���^%-����������^��s�n/���.�$��b��%lG�?)sOh�*4�M|�N��#�KXJ\�8X�0��5��Ѕ=�{�]���"��nfJ4��� ��L�(��#D��9Hug���@(���jׯ녔�#q��v��HhM9n`i�����n����Oi�n�w��'ʛa�}3n��N" M(��3��6�L� =�P��9���n��n{�?�7�Ȓ�e�C���c���i���E:b���)�[�m[qVE�����cjd7�G4��?g�v����u��g�E�ƔV�A���>0���oT�=�_��|bc��@���&�ѹÍ)"N������7S�n:�;��M�ͯ�mndpWt�h���]f]�����
2�?W�^g��øT1V��τj��;��Hn
��Z�P�&��ݦ3�p�8��t2�5��M�haޅu�Rj��5Hy���.��^������h/��Q<�<��\�ԓ�D~�La�N�F�� �������vmK%����-mȞ�ŷ����8��^��GN�2ρO�2wV�O�4�qFH!]^�
@�83�@)�G8��8�K�9�̦��s�ӓc,�_h
Y&���P�=L���um�ZQ�lo79��|I�||!�QZ�T�9�,4�5јVl|��T�y&I=��|1k�%�ل0S�"c��~�+Ľ����|]@��+�N�ã�~�ӄh'����	{/�.���|tĎ<zJ��J�m^�R=���e�Q���z�fg�Bգ�:l���X@-��JP�t.�*>�8�����}��K�D�0�,m_��"����l ���9?|�'�9)�%.R?���˙�W0�P2 cb�%�dm0b��9�l���O��@�,L��%4Ɏ���J����\7�E�=(`v���lP��Wu�2�S�Y�Ğ�lֵ�8���:x�z������*��S<� ڱ��agb���Jv8��s��4��Q���6?"d].���F�����С�|�[�)��H ����r�����2D�>�FѰ���KU^��I��h_QRE�9oO��8:o�*l��ͭ�-.�w���9c@����RL,��.d��$h��J�X�na8�1�Z�9v0�^ى�?�T�;F[jc�l�i0q	��(4�3����ߣӸ}�J�y1>���W��.�����	�#^�����똉J5����&�4`���~�e<@[5PE:�	�^ǫ�~ŕ�c�?E���p'T����_Z�t�@��5(e�٬��JW�1pg���%�G�}h�-U�X���af��q�b���<�-���[�=$�
�,�����+��+�a��q��ޏ�g�;	�;&��d�_p�4tx���F���2ܘ]ʫL����}�wN�<Ԋ�]t6[y��Ȑ��9R>`�����7��H�d-����T6TǀҾ`�&�����|UKsy�7}�I�7����Y|5�{��9a�x�p���*ineu���׶1������#jT�������*~7~j���t>I���� Q��j���7��ō9J�u>"D
͇����0��� W����[*��߈B�+ ΢�hDx|��h�b/ڑH:�� �nCC( ]���8_A:sGH���q���X���l�Xo�����n�&�m��iL��ٺ1��'-"`.,�c!���D�w�����J�����D��ZE���(��N�*��Ǡ�,)GE��}��{/@�/x�\u��,-b�0�G��_�+�%��]�\7��a,<��e\�-�n����խ���o@�����J�滋H�"�	JD�M2��s��Jx��t�а�]�����$a����-֚R2ʲ��Ώm��i���-p�Y����O��24k���T)�5�U��L�^��-����E[/�W�&��T~�xI]�p7)Y�GBѲ(�o��)�I���^;U�[<��7���P�V?�Ŋ��%�i&�թ���Q��L[��d'���؜|�3�&�=�*�XMp�?;J�Mz�x�m�2��(cuz�جG#�@��f�R�\�%�қ+���-!��[��0�֎�y=y�j�=����>�;y|�v+���-v��{i9���j(�v9Trs�->v���V��q$�\���l�s1����IǇv��0s+�ϮW��S��R^�(Ix��L��m~㟹�%Ć�q�GH'�|0�6O�.��>�e%w
f2�*��K�X*��̮D,Q}��~V�5�����'��2TR���v!J��w�������7:�'=!e^�>^!}|�{�9W����JMa?nJS���P���1�l�s����wKo��UZG�G�=����\[l.-�7��M�q�e�xjj�o� �CiV҄<7�����ќ�K�,Z4K��K�ݶ���ވ�:Z�oNbS�^��#��-[q"�N<i�!b�UQ$���\c�۟�Cs�W!x(��G��U�)a2v��5�cԊ�c�6�I� O9�\�]�QEk��2'.�|��u��wP6a$ƅ8�EH�|^�f���_�g'���ie-��FTWĶ�_��Q��Ir;#�;1�~{A�6)H��%���/�bb9Iϙc�W��1_m*W0��a�&��t��S����Ҭ.C�6��)��oQ��+`�CDp�Np�c��̘�3�tI�gO\}�����q�{��l�]V����%sb��t04�X,
�&�,��ف�/&�i��e �f\�1"sЖ�Z��*l��-[��[�a���E���:�] gr'P��7":VD����?'��;c7<?�k��H�z����iP�J�(u+w.�5�w�6|���@��S_]���	�~�^�o���Ϛv#�kxk������%��A���ҳ�X�ɉ�kK�uGE0�U��~ǧIߚk�tU경����hh�l�a���B��sM�s�rp�e����� ����	D6�;|�yt�l�X��9�ǃ�dT��H1
Tk���F��m��	#{b�#�E9L�a���'����D�:��S,9קϱv�$K�|�V�q !�J�sN��S��%aD)!� B$-�|c�f�'��"x����d�y�\���#Y�����&{�*ӓi���wֆ��\��p	1,��Ѩ~��*n���ЛX�i��[��<ZD��g��iU�-��V�n�Z((Q�A�I�ۦ)i��Sk�N u�F�L�1���
��Tl��i{�|������Y!�;�7)��ӱҳ��4�S�(�+M�Nm-��*��_!�r�z�B�[y�C�2�\��{�#nM�qIv�1	��c����V��b�W�h�&�H-O⤯�3�N����d�PA����+��g���'</������B�P$-�̼�`�[B�0f~O�z�X��;=vKs���k��&�������A֕��*߻�;3�࿺?B�q:���i3��;)@�S�(��쀌�I%҉CE-W/U�����9L�=�'��pY-�����X�uQ$ѩU���E/�DQq�fW�M�m>b���)Jmgs?@��A-�o��
���l�j*�*]>�$eǂlu�ٵ��5�Z�e�n� �"����+{9F!��1g�{�F��
U��`��)�'��%M��#\�sk`�SĮ��}3���1{��&�^�`'y�J^MY��?
$G
�$�'�"b���ha��o�}=W���`�/޸�ӟ<Ae���me�����x$��h	h}m�\�z�;���u�nBCs��9�ޜ�6nU��)8U?�,f݋%���I����Q�8�y$�"i`�^ұ0��뚧^������Wpc�l��5#�&�6B���fղps���qpi�Y��pv���um	�MRF�*P��#�,!��L��GD �	�2�X��e��������o��"�_��J.��Ԓ�d9�I����B!4��qw;����o��ar��($�ĥ���LG��f��UJ�L��E���f�c��,���YrtZڮ_����F��^���B�)pw^�w��}G,:��PC�����m�P�rY�_:�%��*�Tz��e���R1
�R&�c&#�&
Pj7J|�=�,�ӛ����Xy��)3Hb�7d-߽JĹ:�ut��D���4��~��w3��[浻���3�$��bY�ܟ���H*�y���cdKS0~c��@v3��Z��d0p@`g�p�c�#qDSB;����Jk���K������ލĪIO��+�[��M�����E�=5]L�qO�f����v&���,��\&�����&^��"wk_�6/�����'��ݕWh����F�9ոq��qL�+���ܨy�ti���]�ᢐ�ow�2Q�}���t�襏�T�,��ދ"rz���g��{���B�΃�+C�5�,y���k0@0$.
��b�;�laS�M��//�|S]��&V���-�\	�
Ib��Q���"�wg|��x�z���H�w�Υ��;��KiN����������	��-���?���\,�č"j{sS-͝{���һc��q�� �)f��']��-g����(�O ��S/�f$»S,g	������FN���j���u���9W�7� �=hHͤǯ���m�� p�}���`B��W�'����b�t�_>�_�D!�Q����4��νkzI-�L��#�Z~�;)���q�
=��P���%N~R�3J�MU��٦��`q����j�<`
�M&�ȃD���Sk����"q���f���i��tv���s�(0ahG�,����1/�[�����:R�"�-�ʢזk/M�k�߸�ܭ�G�M���+O�3���$�zЕ�{a0�+9E�ύ%B>�~���..�B�%`/:A���M��+O��[5~�[�3��_�����BvOe��e��K"�"m��D⿳甏����5j��g�yƆbu{�����Z�X�=�X$}\�.�SQ-�����/7E���豨5�Y�%g`<�~�y��y��_"�k�P�<�@�p{<�'�m��(�����T��m؈!*6��1�s��U�Gߑ�{�������W�	�qDTf�,�eu�@�f�������R\�{<l�1�<�W}FN@N���D;x��b
���vޘ@#�֞G�s��p%��B�׏�uW7��B�����*�ƭ��KC�zeGТ�Ұ���۩�\�A�E&�)_2C0dKj�3��<��*Mʛ�2ul����gJ&��b���o��֩��:�.x��!rq��:?�+��ä��\̔��ܯvɒN]��Lǝ����9Y  Z1Ls*2�m�)�J�{7�|����~����f#��A}�������nh葅*:<�Q<�g����3��j�v�0�ߞ���_-o������t1��P5fW�Q#08�y�ں�����'�����b%|�dz���-]���A��ҳSgɪ���x��G����]�=��>#�n������z�Y�$�$f2jYؼdTk�j�Ȩۺ�>��H��Y�z}�'cv��S���Cbr�0c]��zb�c�S{}�Jq��R���8s~'�rg���z�_B�_&eϚ(�&����k�Z(�'�L���e�yND��r#sf"!���.9´�#������N�l�W��0�>j*Z̙��l���|$c��.��<	#�K�t�%�]�w�W��d6\���E�!h��cQ���+TǱ��J��)g*�AO#߫)@�F����#j��Dv��8�1�#�������
���������q ���C���{� �Ĝ���mT��N)�bN� � u��T$h�TA��!�O0�>;
m�l=�+9o��i	$ĺ���L�9X��]C���!#��U�Ow`���_��u�1I<B�G'h����j��ȇ����������;�y�/�c��M4����D���Wr-g���TOT��x�Wqɑ��	{O(A��a3�\�to���F�l�d�)`�/���9$�1Sy � mؾ4iYzѼ� 2�N-U ��v
�� ���O���w�G��O:,\��z�|���������=�U��W�K�?^�N�9��&���
̹��D%�.ѐ����-���r/��8��0R�e�����3�t=}98)�PY]tb�1��K�U���&�-F��:YAyg&���'�?_Y�[�C2-;:$K�J)~`�SN��8n���Mi	���%	cA�����
�y���?W�B�e>Uf�t�({�����d_�\ŬI+#+1;��fD6��Y�Vj#��Y�L,Cf��/YCoȃ��P�5�AJď���<a�X�����Ȭ���SN�L��z�1r��&�p�3d.dm�;�e�_z)���?���<�S�嗕�b�/^��A�geM�R$D����1�Ox�!��3�#pKv����aT&;��U�c)޿��8/�����%%�h��|�j�i"��@#����槟�ŭ�
	ꏜ�^{BHaRԸ��r�ɼ�{qq��hF��/r>��~���.��G��f�G���L�LYk1�qY��g�J�LS��u��P�!pL��_{�Ĺ�P�ٵx����nL�n#�z?��q�[/�Z���*�����"�c�����e�]�{�2�ȂPəE0����,5/ϲa��җڌ8U�L��6��W�2eM����pG�3#�5�|X��+���"O#DôZ��5��pk�(�0�e�����0��M&(j�J��䪟�k?�����dْ�ēz����~QT�͇�������P�]R)�;�P.�nν�ϻ.��Τ�{���0v���B����¦�m�a;#��T��=���͗�&+���ݷ���w�8Ʋ�<<מ��41+��+{)��z*~��ASJ2䍄KV���JJ��&m*�9�ЂT
8  U��ͩAEh|�e�Pj>����OW��9�T�}@�\��9,�t40ș�}g~�p�K��*hV�)�$)���>>��DC���E�@�x�gE��1�X��s���i�E��ؔ�6˻�Iv�l&��r�����& ���筇j�k5�Ъ':����-��o�P�g�����c���e:/;Cr<�#'����w�=��H��0�L�hJ�~ ~���Qo�)�Ջ؁����?oMtDx�1���g..�;G�z1�R*>x;�u}�>����歐"ah��[��x%@a����|�������(Ll ���/���1izI�!�4�:(���v0�h�����ï;wU��{�6|���{�Qq׫X�q��Z�m3M��1k������P[p>�����V'hP��(p5��Q���,�� %��+����&eg^��������L�Gw���X\
��)�q��r�O�$Vo�������'�4�7˂e_�ּ�_��2k��-�1"D\�)���
��X���aq+m�(��u+]���G1�*g[�k5W��^�������;X�ͭ\	I�@"d#Z��4��K3��
��Q���U./��Iw�e|z�eSl;\������x�:K���J~Td��>���r�uPuh��ד�_1�#�ƨ����kbJ���p���" ��t�PW���u*�&�I��4���E~z?'Kǉ+_>�߭x�P)R$b<� I�
Il�´]�������p�:�[���������PM9*a;����z�PRD��>�਀����=���p\��v���N^
LxLx,5�����G ?=?1��$SK� �ګ]��*F�l����ϊ����ˡ���]���������~9o!X���Je���-��M40ޑ��D~  �VLPL؊���WH��i�F��hX�O�=�K/ �A�%��Ȫz6^�R��q`0�bd��ۥ��x��b� ��Q���<�ta�N�qX���H<�E�-�t��L������F�J�}�<�0���%�v�8��v<ѩ�"��eZ���@C.O�������`6d�[�� ( .�����F��%��'ؒ����Y��cs�m#EH�/�^G��kik���ʡV�1HmZ2����k�����^9��x1�"�˺�~���V�Um��ڢfG�
�A��(�D�__B]�U��u� X/��������nb̌��H�T�P4�+Ѽɔ
�e����fz�-C�K��WSx�qh�儚��m��0�\#c�&:cZav���ƑL�eX��R�_8�Zk(�(�MŪ��6�#�q-��~�����	��Z���c�MA�y�E3����E�V,[��(s_Sf�ik�2�>��SA����cg���E���ݍIU4������e���\� ��_�Ѡ3��������%S��T<�(A��e�����rG����J����i��[f�v�0:�D�kE2���m�F�B�m�K� K����B�x��x��@�7�g���ŀh �2��πx�`9b�	3$3#!A�xi���Q�f�'�@r%����u�#Z�cƔSH�n�"����#{��O��CVB)=`d��H�U
���d�����&i�����W��F�Hhp���)}�+���B����9J�������Y�>z$�;���IH�(��tc���^ϊ(��k�A�[5��:�b��)������ ��mPI�g!����i�	� Ɓﭡuud7X����Q�Q6l���� &P0D��k�1Q�1�ݠ��#U���/��	W�4�~���|����������#0��]I}���~22�8ZN2��2#q��|�P9	��=
�H/����C]s���O��WD�;��B��f#�ϻy�ʳ�r?\�ӻx�y���&���pX�#���ٮl/�cW�O�?xF�֎�֮l�+I�+ǁ5l�~C��|׆�zX�jF�CՅ���?r�?��$�%��[%�ȋ@�zbB^�L�����(�$��͛ޢݪw�@�:߅��Txa�p�����p�a�XwJ�R�':��!����Sb����P�|h/n�?)�5Cd�,��Mb�ߠ}fŊ,�W���H�|+�0�^�:�;G������Waq�~�_��/4)��E���Ç�Aq��5+Uho33��$lt����S��|qFJ������9����[O�g
T}��8h��Q9�P�/Q!�Z�י,ĥ�߆��A���q��9��cbs��#U�h"���D�5�����季47i�Pf��ry�L��-���y��u�gcN ��R-��<2�����-+�K.
�������m�p48(��bwkw��/E
�b�+�p�tL����,uP�@�G}�LfE�"(ѽ��9dm�7;�s=�bD?�nD��f���6�L~j��n���{�׫᧸�.�uю�`�xΨ���`oE[$�����v�ؓ���r��^�ʙ����<ݩ�1X�ʐۇ�ё1��a��M�r�)��=�7���eOj�_�n�[qVcR���k�"�'RS͆^t�q���6������F5��Ϯ���z�X���f��l���e�f�:�>|<�?��{�|��k
 ]#�a9��F����GBKb+��h��L9��x��K�Cػ�������2�<8Ć��y��u�^�~�7���5q�@w�G�d����;o���oy�K.��1�}X��QTh��Jܲ���j�H�M���7���-$|��\>O]��(���ܽ�7�2;����y�<>(m�w��l�� &��X��V�$�"i�c��	��K�Pt8��5��5���"!s���Aqpb`�}r��;@���Y@����T�P��ϡ�j`[C�_R~�4aG܃���n$�/��������/U����W�߆=%�-�B>O]�����<ޠ0�[�.X$z�`���>�XXx�Do���0����sx��T����zO��f!�/�VoC�QZ'>��5�;��p�����٠3*L���Y�Oɛ�/h=�(b�GHl"0�,x�,�	$o7�AHm��,kM9Tcc'6*�V��Q����LM��u�X���t�p1��x��s���"�Q�k#��� tRI��.5=��D���"*�G���n�ϣ�DC2���WR�k%R9A"��w��

&TM�0���kZ�g�#Cm0<ZJ9�䢳�j� �:1����;���n��GJ톌�hS�	A��/�(i!Ԭj
Ʒ�XQ�n��y������\	�"rҐ�����U�l�@@�耔?�U���$�����?뚌K��,��7��#�<Ba�M���c�������	v�j��Bl�����������v%5<b=r�j����ك��3�Ա@�b������inQ"a#נ�a�$��.\_8b�n0��ē��+� ����"�Y&�
V
�n�x�]`��?-�@-b০ޭ௠�h��s�&Ip�?MP�YU��_�U�>�D�W�'�^[͸��J�7�� �\B�!�����48�9��̥�F�:f	t��vZ�]�o��q�a
������՚ax2����԰n}X���Y��^�A���&5�M�
�X�O=^5��ضN���*W� e�����4u��Ll����F����n�i���h������0[H�]	?G����@.j�Ttàı�+d��rO��� �c�-��OF�+�T��ϣ�9X�
3��Թ6J�軱�i&C�G�Eώݘ��g��I��\J+(�z5l�s¹3q���2S�b����ҹ;\���F5�:oF���&��0��!rWf��5��Ħ+J3� "�{��P���r�|�Ⱥ��B���yz��%���LF���o�`��M�T͢DE�zp%�
x��[~����$��i\f��1�ǖ!B+!|��_�(-��.a�O�~҂I'��Q+gWF[�ȉ8h���~��{��;-���9=ul���W��N�v+�>�z���*�R9AZ�=��x�'����*{�[��k�䷴�� �bu!sZUC-�a��g:p�:�+T������=�Q�v�B��@�S�t��R�ڄF��^橜�e(��݂)��1�����t׮qiΟUmڷX���=�Nz�$H�9t���1X�B�X>�P}�?��d\��	ʎy��xZA���1M�%��U)�ک�[�U섎�@gB�Y(d�7}�����[Hn��lPQ��2vvĘx��&�i��{+�X�"�'�����=2
�i�`�U,b�gf����G�l��"�#����xI�;��鈸��A�,5;@F����*�P�m��&���������V�k~��K�- ��p���x�n:�>t)� x��M3�)�M�l8�-����KG����8�`UI?���`s�F�p�2�}Z�����O�Kc�f�
�!pӪD%���׷�H�
�8}�Q/�`��>z;C���49fjEPo���X�Dr��;�5���^�[� A67�>X�R�ny�7i<��PI˞S��xMx��n�X�_��O4�d׽�0[Pr�eT��⽬�k3<nvGV�P�^.�/{5^�r[f̉�6�y��y��E�YE�G���*���Ur��%���`��Y
�Ʃ�@�����F1n5�}�z]��<.�W��D,J�d銛a݇�Toud���:D��Y�$��6�+i*$�C��`�S�ws�c'�]!L����qZ0<��Ȃ�u�Nw<�����D��Uo9�i��ş"R�!��,;�6�\(Ճ>�X�>�"\祫=�Ǿ2���`����_i��S̹�1� :#��j\�����[�'��f���ن�V㴴"veў135=���	����ɧ��� M��`���c�5|J��i���'E�)27�J�㯐$b�)��B&)U!���f��A�m�4�!b͆�qi��}�����J��9O���n�8��
�tF^PG���x�\�x�[c�v�RP"?SJы"��q�r����$��Y�l�(�-�P�J1��^	CM}h�T0��	�P�Cj]�P���C}a&��l���Rگh�����@H�.ޮ<ֹuSC�˻Y��h�Ш��R���.���=�C�X�;�J%V�ik�W���z�m�z1$ވФF^�7^�'ۂ�1����j�B�tJ`q~g!t )c!�B��|�-�k!�Q��O\�'��72L+�|��[9�VX�7ڤ]<e?K/��@/W�Z ���d_-Du?Z�s�S2�&:�#�$������tJCe��U��M��;��F��x�jdwv��ѐ�8��7�
�����1��9�-����"ɅR���48k�nն-��\d�p�=��zd)�hk����ۧ��+ �mT�v>�w�t��7=z�ʁ� H3���F�K�#L����@l�[Q�����6�2d<���'D�T�F���-mV+�#�&��0K�R���k	׬��P[f�_AnWL�ˑ�U*�u����$�zfz��F�Ah���B�Ǌ7x����ݰ"�ne��u5�B<7�++�����20ŎW�6�<����ܑuk�����\�@�B�)+���k���M���J�\KFg�"T�"�E� h%�#�T�  ����x�B�,\�b(g;���}]�@~ݍa��V���$��]�+9��FM.I���7��3Lp�e��sfn϶���bs�+������X�4�y��� ������8�����"�$�	f��ri�3������MǗ�W*����P��'R�t"V>�!H��.�҃e��8���ܳs1�� �뚋��k�6'}b̧���3�!.ko/DK�[Q#g7��e�
�E	�zzh~�p��7LP���-fv4��?�L������5��zw������Lӂv�~�F�:xe�~��;R�r��|<7Dת.c�~(r�h�r.� 1O�$� 3u�fj����(3m����N�>�l�|o�)]!�K�r��?�F�ڋM�~��u�������K�$��8A���F�ۂB����E����z���%:|���Tcnt�Ve��=�)[�p(���O>2�W���u�m��Nt�>>H����_C
�k�S������I�/��l�4B(������Q�lcNx���#S6A�s�d�m��6j�-�-,�C�7�Mr�x�61/x ��QPR�L�㱥��;�m��(=���
�#���ǥ%Q>���/|��O�,����F����\T��L���k~j���@�����u�.�"	������G���Qͭ��a��:��e���>�6���m�NU�1���a/�����d�-�p�ȟ�t$*x�hgl���{X��[7#�3K�*�~��Y��RN�7*+�	���J����L�������Ȏ�rO>x"�.[M_�	_���/��SD3���/�K�+Q)�РK]���ճʈ� S�K�gf�܀+�D�k�y8x���o@ݬ�	(����|�#� w�8
l>��������3
���f&����Z)�ϲ�"a��V�����' �=��e c�8����]������0�O�h��y�"�������W3M�A��\0)k�ET3�q�0���>ҳ�=FY~>�����:9�_t] �;�ne��O��/�X��R: ����uЛ�Б��ۨ
��na��y�&�{�RO�]��p�>��[
�R>�����I�d:�H�N�1�ż��՚ghM��h��_""���<��lHaoh�/RW�;%��Q���g�J�r�
�F6�1�9x�m�����+���0ww	��������5��;!�����n�/�n�{ﮮj�v�gG���z��y�?(訩P]�Se�[�P�x����8�>��R
e��c^MI��T���7�#�ʌt4���h�#U��NKv%�9L�U�.��9�U����6��V�B\�ِ��H��b��}����"y)��tϢ����m�[��^L~ng�p���;D��|�fYg�՚�Z; -<O2.���{�;�� >���Sr�$f�X�db�ߧ��sP4�AF(8EH�v�ӧ�%��&T*T�u㋐R�tI�=�����U�|L�f��]xL�.mL){Bh���$�-)�{���ǩ�M�++�M��d��G��ik����@%߬5B���Tk��#l��$
y��f� �����*~�~	�h�*=Y��fܢٴg���ǐy�Cذ�	gT�F������~*gC 54�C�/��$6���y3�^yG���>L��C_���W#2�#���8"�V����z��hm&7��sD����T� �e��Js�@��OC�ov�$t�)� ��*�@�Xտ�$�����%�Ù	`<g,Ql,�����S�2h�U�|���e��Z2]C;���s��N�7ҕc�~�Q:B�$C[���F�dn@L����X��/��;i����%��~l�*���L�G����k�
ޕ�F'�)�1cD�9'Ș���f$���F��ؤ�W�_�c�>oz�$񾅴�E��0�����*�7Su���G�]��3(�U
��'�@x�*-�^чY�ʎg�!�Rѹ|gCĞ8�̈ޣA�
����o�J�%�)~�R�x�%I/��̷�I1C<��20�kg��Ӵ�l��i�d��CM�3�_�D�<�|e��O�kII�_%�j�^7���L��ߐ7�T����B�є�D�C�|�`(����e�B��8�-���F�G>��2�E�	���K���C
�t���$C��;�5�uQ�!.rX�W}�҃�YU��8ԳZ�&�{��ږ��x�v�Nɬ�;S@�G�P���%���d���x�|g�}�t�a�OWC!�R���~V+�P����o�HkbX-\5��՘�H4�%e񵓥����~�����/nO�[f9�n���	�,	�x��r��Qgְ	�(�pH��$�5n�>(�}��'7Ϭ�{q~�솳Xı���!�\�����.$h>� X��S;ђ�o�~����a:��c��pzT��榳����\|U0L;���L�pK��%���s��.���v:k6�ٱ�R���T���3���Lsь���K�o�9�����s7�\~�C�f�*�h"m�QQFK1����V�u�0�,�#��Nvc}���xC�9P��C�_8����^�&<`L��E5�ٽ}�޾%�_zJ��dP�7��C�U{s�SP� -�e�l�hG��p�T-�Q��:��tw��d�f��j�\�"L�����'�е�d�з���J�P�B-�Y�Uh~-�� ?nrN\���8�u3�7�z�^jԷ?�_i�uJ�~ū�)�����nL�]����`�:`��|�թ��+�l����+��k��'�R�h.��;���**#�0��,�D���78�)��%F���EV�*����C5@����P]s���	I��Q���o�i!=�A3p�h��I���
e�߰R�y�oR���KF�^R���1�����y���� ۛ�I�(Π�W���8�#m)K����ۃ���x���=-������nS�8��ܟZ�&�D��4{d����;:?d�T��z�����k��I��Z�����an:��ԌP�����7�g�c�fE�5�[���M#G��D�<U�����S��0D��ԁw��+TDi���)6;CF��5y&Fzc	2�sr1R�p&�����鮆R60��T��s��\����|�~��������U��cs�ϝ�>]��ރ=.�i�g	���n�x_���BI�L���IoƔ�C�^������RVDY���ܞ�����5�^�
ˏT�|��5��T
�Ԃ���TTV��t�G�)���6>e�|g���	I8�Fm���S���^[�n2@��ݎ���R/O�+$��nn�-�@,	�����}���`n���4F߅Rw�� |�� ���X%�R~�T%nLO6	��4�df�w��[��,!�[Du��UŬn��!-�����u�N��ςz�m��\9����wh�`i���,�Ҁ[jz�3h�rLJ�0vۄ����[h�+��FE��}A{Rp;����~f<t��	��Qmk�Ty��	����ַ=��AcB�%�#�c�8
��?�m�v�	�N�VT�3��C��}��Yẜ} 
��(J 0�C$�V��+	\�w�%�'T����l<��m��G�#�Y�.#>a�X5��q$��E�����D���`�{+�#,��:yi�8�=)��嬿V޺~��m�������:b�E�$�*�Hۆw�Z)�n��t��� �p�!��q�B�"��椴�X�Bx/Sx#��4x���4������*�ɟ�`@;�$� �zU��M�(rtd
��u}��d��/�J�3Oy��T��s����l>|p*䣆j2E����"p�N$��H\h��F��?֯,ܘ��P���+R��*w�P%��o�I�i,׎��a�ƫ�������$	�����.�RǦ���>���,�D҄&���G��k���w #�
á|�6�µ� |R�._@ _�FV�>>W#/������_B>n�S���J*fk$p���|�K�j(��8�Xǖa�x��q��eG1}�3
�//I�:;��	\����8Zr�����rE/�t!@fu �^������?-�q�I�F��s
[~�����CS,&�����&�0fp���ٯz��H������=o�;��vgUř�WĂh�@�5q޻�0j�d`�O���ձu1����e�y��!��dZ��`~Ÿ����C'�MR�t`��#h�#.G����v����*?/�����^�
�N�^8��O�2������&��6d ��w�m�LK�c����pS��Z�ڨՌ+KP�`p���=�ТY ���1W��9V��?\�����\�R�\�V�s���-��av:}�*�����[�s9����EQ֏>�/�	?��f�̻[��	�!%MW��xm�d"�Q�SJ��� i(�A��~�Oo���#s�&A���|�ЁDϥs0>}��r!�*��D4˗5(W��|��W>�G�ợ4��f4/��e�s��l�I��H���]�t,ymo�~Տ�Nr��t�=�Z`n8�4���k�L��Y����������{vN8?�0�z"�G�W���`<����5���>�,.��(d[3B�:K �;E���`C��hO��,�$�J��"%���X��q��"�.v1���iP���Oc|�C���.�+�m�c��|ٰ`k��ƈ�k$�� tC�e6|nի��4L�'>�t�e�-�$z~���;���+�ֽ��Rm���ZZ�w ���JM`��&�Q��h@�U)%���yj��0�G��n��eo�~��m qE;C�;# ���/���B=�,"�
'@�%��G@{���:�J�:7��E��=���Ly��s�ߏ��\!�~sv����F@"թ���5���"�I�|����n)�&�ϡ���s��9Tb��OPվ�s��"s^�5�%�A����D��p�FY��O���Ѱ2�rI���h>������s���]o�TR�߽�u��z��������t���"��ڱ����?�p�a�fT���=�r�&Y�ݑ!����S�G���bw���k���(o��x
�d<�+&m�D�"�ȰPK�{��p��ѡ��M��S@�q}�=h�ׄ�y>L�����깴u����A*W����0K�M?�/ j��m��{T���>xVf}m���rh���\��\�U��pl�XE.�l�H6�Js_����>������8���iX6 -z�˴��n����MH7b�����7[8��M���K"�`����d is0I�hQ-����,؋�Z�:c�ݛbqk� ��{�|�����e�������M.s�����	��3�ϥ�� 	hW��9с ��k�=�|8����ȡ�X���Ĉ�s��wmQ�&R���[�^t��7��m�%�u>-iӌ��V?�`�����c���ܴ��x���OtZ�@n6ȁ��o���ra$����\|���)���s@����)����/�$�3�*	��f�9��uz��
����n(WG
0Fj}��[@<&���q��lq�L��[{I	�ޝ+���w<�����KK�Ʌʱ�ރ����E�7�ű�&	���%��-lHZ<����t������PX�mݤ�����d$D}K��5�%�+�L����Wk��mG� ���]�)��G������m��n6�L�f��[IX�}T	�]Hl��(S�����:=gư��I��۸�N�'��]�!e�pG=��Iq]����C��bܓ��U�����2����+m��{�`jq�h�FYv��Ajn.|��B�"0^�.�!;�<)��\3ˀ���.Kjr"�gCu�md;]i4m�?!/�ܾ�$��N7�X��1���CDOBM�8k�A�e2-6k��&�{˓��Om��My�ywvv�����H�|�)��TgF%�'��=k��=��ïA�`�KQ�ZT7q\2vk��U[�!��7O?��]"��a�n-��:�#R��������)�x0�3_f��
�D
��a��NoM����wx^���S1� �߲�.9��_��MK�v�aJ�x��d�
�,Y�X�ȫ��N�=�]�7E�3�E�l}J\MCV�#�b�>��=�CM7���c���t��A#/3W
����M0�[VP.�{����9�� ���Ck�O���h������OvEߘ�̷��&�I����E4WcY+���s��.7]>t<N@ J���g�z���Fce���)||�.��Q�5�,��*��$�C�v�Z 範g��d�ໂ�z�-Ԯ�#�a�T,�h�[�*K�P=��C<o����u��B,��	�N�����k��6�z8z�y�L�ʏ��ټ��S��('u������hؓJ�oع�ȅ!ӑ$�O��JM��P��!�Y3��Ƚ�3����ɟ{�,9�{��Z�����������d���:�Rˠ��%�e�bg��uD\𖾇��gf��8���
�[qI��d؜�P�.����4'H��P.�Q%|t?��"�w;��Ҽ5�D�l�&�Sh�J��Q��F��~L?�ȉm�s!�A��Z)�޹E��{ۇ�G���8������{���J�� ���E�#�������Rb+�4`L6�G�|��F�K?��r�g��IWйH^�q-Mn�s=u�۔�d���3�&P)�t����O������x����I�g%~6���Y=������5�9z1>b��O�G�w?Q�|�LP��l��U֢|��#Tc#N:#C�|�v�\>>�Dk�W_7�&P�+����^�>y�ݳ���W'�Dfh@5�³mнVe����[K��B�6���]���u�JJ�B�:9e�q7����/��3*�r���8��B�GjwP�G�U�)��ſ,��:W�;��qaݩ8`�������%WQp�])���Hʼ���G:� ���ViN��S�D+��b�6�?�a���3?]*�r>h��<��������݁nX��"r�*���Ɩ��˕|� Z�A o:�?�x����>2�~���l�#ξ3y(��3�V��� �Ԣ�
���7�Ᏹ̙8��L����徾��q�U�s>�p-�٥{,�˔x��g�Z���]բ���/���,���՝���qsu��`BHþ����5�[�ԅ�������|�A$�a6�$fB���Q���5�x;�F��G���c�B�
��6";ĺ���
��oW/h�3�x�K`����\c�Bם�ul�s�)﫠et���[�U䌄������&�܌n̯g���(`�E��rqqI%ѵ�n��G��$p������Ͷԩ�\ �e���R74990�؂;�+ֺ�����W�3h��էBO;/Jb��<��������[�j���刍3�cM���B���⺫�Z�|�s�7��}�[���Sjf!���sy��`\X�ɾ�~^�k�VeI;5�=R%���V �g�#Tk���C/��i��!KL6����ˤ�h-�)cv�5�g�QB9uz�>�0D4к������U����u�aA�ns�KE���Y-���:P�I];�����@���/t�=.�r�6�ʧlj/}�'_1�
���P��7� ���S�l�����r���$!d��tpXr"�Z]�]��^N�(@���9��t[�Qvz@��fD|���$����Q��{`Ne��k^l���`YJ�=s�%oqg����������៾��;��^s��ȥϴL;�e1L��(�1|��{���w9!n'h��'�]3h�]���
�
:NЋ������|�A��wd�(��T9�c�s��*�M�sd�����7�To�a�.Au���H�gZ <]��ĭqǍ���C+����廁ҷ?�ڪ���&�bp�)~��2�/ʸ��45�e�Ҩe�h����3߹�<O�`�F��ߑU��0Կ�z�q�I�ND��w�xq����PP4�d�n�]�<,���xI�:)I�ވt�|�o�7P��?H���cסMA�t%C*U&�m�����J�i�ONI���9�%�S�����y�H�֮v�IU����bEq'��<�"CKh�,��IM�<��NȆ�h1@p�8�D��t& tlg=<�X��ИKԡC��;���{p��!����Gڎ�������o������3��j+B�����۰�f3snbxU�|����3p���}�
ɓ%�I��n�N������M�&�8�ZP��eԸeذylKM��.B�"@���*'��M�
��=�CR��&�C��CY��5��M�n�
�.}� T�<!��s��(�G�f8�+���S�'e~���$�-j�yk4}s(�
��F�:���{�!ʫ+�D*6g����PTs1�5��l�uR�&O������d5�9�И�=rũɱg�)B���ir�{8#q�����3CX�{�f��M%�x`�'�BP� �K���lI�����9����_���9� SG�;���0O�<�z>�f� �]������D
�f+�����wEy�ǔ���-��'0��w���,�ʌ޿1�ډ�� ��d�	L��䧘],��|�'P����S)Q�;mTq�О�H��.�Y������Y�/�������� òu���j�b!P�4,�6c<ܩIs�6����x�ݹ1��ڎ��J�,� ��%���18t��E�&l�4<E����F�[�5^ٟmvf�2��˷p� � ���<��P靯���˸dG�>\w,�F������W�^E���Jx;��=���/&u�7u��r���A���|���ɼ�0��1���r4<�w����ƪ���YE����z��S}HYY �҈T��Z���/�:�E̰qI����:���h��;��OƗi��Y9t�w_ �|U����x�]�;�Q��<�?��<a�C�-����Ҟ���E�X�|Ę�{�rL����ƽ�����'��$v�I���l%!JU��G,F.�"�|P��i7<���G91�����-|Q��:�W����)`��2��ǔ������^�t�O+�X���xzY��1ҋ$�|ْ|�>3m��0����/��^��6	�(��V6A����z���������g�v0xY�X8
Z$X���t���Di�1�.�2�[ק�ݧlT��\���G;�s$ǋ�S	Q��2��H�	���Y΢e��}W=U�ߓĹ�	�oN4+��=Ĕ��}�Y��J�T궴%�3���x��t���]�27OQ�>�*�7�`0)ǽ���Jo:s���K��@��W�f�x��y�z90$�����ǿ�Ym�Z
e~�§�$�l$��\�
�lb�o-�l;w]>D�a&iMM��r�^�l^�	N���>.5�|H��o�.�� ѥ�}*����.������ɚ���-�o�]��&6�`�1��-��P]��k��.s�������P<�
���~��:O�6������.�<���?8�@W��@dg���n�F�{vl�b�d(�6l[�h}�8#�O@K��� e�'���$����-��M�(nv�b�"���R�[�~���gCSQ�Qsr��� QpL�S*H"�5�g�)����~����wlHO0�1�yZ��"F���@�'�o��9�]�o��Ij<�@?�Xyd�A�z�HF����C�����V�"�tч�ͬ���)s�n�g��6@9���}����1��	(�-] /�Nk
��߯n�?�!��8QL���\�dG��xx�z;��L{��aS$���|�2_֛޽��N_��/��5�o|=^7iz�8_1����f� w�#4��x39���z�)a�ڿ�$�t��wH��ƈ�7*�V�(�.Nn����Q���b[���ӿ�w"��.�vP�w���]���2� �v���\�V-*,e�=���]�s� ��8��;�#|�fߢ��t��;N[�C�ݐ�ܠ0?`�Ƌ0�wQ����"�M�<K~ޝ�}��"kn:�*-�'�����Z��5�����/���;�S��u�v\�my�!h���H�Ò?S��m��
1�����-%��v��>���0������q��֖0�Y�X.��f�{���N�%�@���"0n��_��$�V7�>��&����u3P�&�w9�I9�{�c\>�s��4O�·C��W��Fe�U!�V����Ȫ�av���GHN��T~�����g�����R��V��� ﯚN֝�v�7�</�=#�!$�[X���?�����ޘ�<`CJ��ú#�31Z�nD4�a���1�����*h�>^O��כ���K��^�V~�;�0�c 1`�w�Phi�%԰�V絹풦�����K��E�1�H�����W���nHJFUTk����0t}�Jn�EѸ�U��)�M4>�x@{` g4��%��xC����R��R��d!�t��c��d��["ᷱ�HK�޴ o�KM�uqK�� ������b��)�5��f{yK�b�K�g�j�����^��A�c��ȍ�C� H@���F���jѡ�VԀ��R���_����]�U�l��)��������dN�|���C�?�+G��9�W��61�jn�����V1�Z�G�ձ���hE	>C�ӫ�e2N���rw�o��s�RVQO���z�'w�]���Bk�{�?��=�Q=;����?��(Д7]n=H%�9ONϒ2��a�� �b� ��8Zi�p��^�v����#m�8�E.m)�Q�b2g��~S����>��evp�A_Z����r)Ó�?3z6�me���O��z��xn0|�*dE߇����0�r_��%�z<����#u!�~�;ۜ^�JF��X�"ҩ�v��ޣda��]��l����8t���F"�V�Zl�M;C&�9���{E���O��vjs����2L � ��7�v<��>��e��������9ݥ��+q&\�����V���7r�%�-�ѥ����ԉ��X�i���?Ü��.K�����J���ѯ\�Z4U���l�$P ֳ��O�O2�#�r9۬f�6��;>�xH=j�DR�)�h}MZ��C^�u�k�8��,l�����;Sߌ�����{�䟋EK�,�[	OSaGN_������TR�����S�@��6��Ow{��
��<�%c�<ޕ��|M;p#Ƥb���#�V� �,����+L�P嫯s��k��1a=,�JNcP>]��\'�.�A1J��u,���������/ˊ��q���o�.*/�co��[�Y�R��-�&�Vq�*h8�dcW����#Y��tX�ۂ�Jo�z��=�0�e
*&�S!�q�����$������k��4=|_��8T�c»����a䤒[W��Th=�}��;a�U$򡚘~N�HtRi�6m��ᬽ^c�z5g'?&f閑�OV���1�� 4mZ�+�2z%#B�BE���%��l���i��6�Iy�"�p!�W�b�J��Sܗ����ܶ6��݄f�i&��aõ��z_Hｰuzz'��k��6�9O�P�t��r%�Qd�|ƒAp����>�M���h��։B T�d�F���{|e�0f�$a��{�i)Rk��R�O�<wsYuC�IY�5P��34E�%X��#��9���^	�a
,s��b(�j%%�:��t���M�e���ݸ���qȕf�
�q�E�銘��~8���c#RcZ����QS1�YC�������W�8l҄gPxD����P2�6�+��voV)Wv�e��6a� �c���ܸ�b�]ƶ��U�þI,��>{{\ӟ�Ԯ¹��1)������oM�g��s�Jn�����^_mE���\L���D�G��s�wQz��8?:����`k��tu�8=!J�
��� b��3���KG��L	�8�z� �PK�t�lC>x�Ɛ�F^j������=�>d�z�B�S�0'�nm�2�+IU�a(�3�|��ͻ%֙�1qj�ƩW=Q�Zҋ%�A���:� p�]�;�v�}	�&��>���u��z��Ֆ{-���醦���Ax��U��_Ȅ\'�V��bu9�w	�Ab�u	�5�SzFT.�Ԅ~s5��l�O��o������,T%��$�Օķ���HA��;l�n����n�(hy3b��q��ﷻ�4���~G��2������ۑC��� �XR��	OC0�/nC$�I��^B��Bp���x1�JBe�So���Nqr 6��>!	O|�|�8����gN cy�<��D��J&�,B�D�iH9��3�%���G�61
'�e�T��
t[	S��D��=����8���N<f4���M�OFI5$mGx��{���R7�³k	�gϗ!W%��#��2C�0z�Zi�v�(y��z��/Wd%��@y��i°ȵ�ߔ��d�/:B0���e,$~�k��p�B�]����Q��Y�?����d����p h$���MSq�W�k�E�/`�;��TH쯂�N�����ǿ����S�Jp����+f=_����ݴ�Fzѝo�������:�)E��LN�&֌��{�n�1��M}����@��*1TƎ�,%���֍�]G?�|��1�p�z�9:��+J�b�Ӗ����G�Jv�f~�I����ټ$�v~ڿ,�"��mjs�����*_��N:��d�1�#?=|{�ڽu�9��e(��A�p����*�ۨ�����a�jv�Q;�.��7�B:�*h�mkO8�)�q��4�r�W����i8 @�	���\���{��yA��M˦�jDz�������1ʿq���=0�A�%%����BkU�����1�B@8z���@ԫQ?]MF��x���),x4�,+s��v�d}��G:�����@?�a/�~-W�OaW����s�����ϳ��$�:���o���h��9����g��&�Na����ho�� �ll�s���	�NO�p*mw�|Q|���`�� ���?z3+G5b�+6`W���y���
h>­N8>K�xJ�yQ`d��#<9�<��,��~��$/�f�b��Ts�P��^_�t�?��R�R�9�VB_�~?'G�(�s��X x��*�v�k�N�>$�[�pQ͚�D���ݪ�
�w�����܈	����품;��]h����N�2R��E^�������'�z�ffL�b��4�k��	�{}���G�rI���"O�lr��]�;��?8<;vߵ�
�Z{�og�˸G� Ѧ��V4���p�y�Ș��_���%����D��������{��2�5��{c=7��u��?9�F���J~8#�4TZ��z��)"x����_%!������aA�*��|"���
8"!��Jv�_�D��t��0���ņ�KК�1�֙z�A\�K�}�7�y��6����@Q�;T2�e��fM�	}7Y	U��UI���� *������BY��`,�L �ɇ&��i�}�e� ciu*!�\D�wԀP܀PT�6��1�'�5S!��x�,�gF"FiL���j<�|>��������N�q�-[^�&]&?R&�&R��N>ܐe܀�m�j~+�W��T�������+C�i3���;���>EقL�}K���p:��.
��K8g~���3�\=�����c��B}�$�5w3�9a���jOtc��p��P���
��s�p?�x�H��$t����k����TB�,��_2:��v�<נ�<��K�q3�見��2S�5H�����ʊzB�`M���v�F��z-�*����zl�u�=�HZM�Y�sc�����%�w]că�pb��D��s0D��`_�����{��W&X�y��n�
pdܑ�me���ٺ�R��Q󦉃��v�D2{xtq�u�L�I:�M�4�ޘ���A:�md=�s��s��Y�Y(nv*�<;��툚y�:T/U>ji����<�\��H>R`T3!��w�!�����d�Eb`dd��V���1f3����JJ������	���D6x����M�eVs''�b7�%��B]&铵$��6�ɓ���� :˺��V%=��)$8�5c��.:paϏ�6�K��:v�GgD��ms��;��|^����>õ^���6^����(�6�������=�������������j�g:�~ȊyDpkӃO�[�]�=X�r`�\��y["�m��zٞ�Y~�s�=�����-,AfTV��ʬx� ��V�5�����\�y~<�!$z)M$���w�hs?:J�h¶c��_LWߒk>�#���ri�<=/�:��OIM���T9O���׼�ZJa�NIH���o��r �}���xy�+�bEDDL�*ۣ�CC�cKɦB_�3�!��m�@6�n%��O*U��U^i)�e�������
�����w�.��HC�%�\�R��!�J]��XZjr*U��&���DK�k����^T'�ν��D.�k^�� �ũ����P�̭s����-��m'-�Eh��JE���B��㢊�G`��;gp������2H&0Pddd$O��\�`��g��[;=���a��]�X��B6f�ɕ�X9�,���B�e�R�]�.��������s�S}��h��#�C����འ�9�������n^^N�A��FT�k�?	���9|���Pbfw�p��4)x�����=��RP��(|Eظ�>%/kf����f,c��J�/����x�D�������l�#��2 ����=V����L�^����\�zNGG<�/�G<�xK9�ŏմ(�Ϣ��ClQ,���n���d.�`��ś�eai��Eް������s�3�=㯵b! �FU�Qn),@ӛ�\�sЍ�턌~�̑ܘ��SnC%���ŋ��j�v�:�`��$�U��-`hE`d<F}��X�y�hEc-hlą�8:9	ݼ��,=H%����z���|A�����!Q}�"A#$$��T{�l�a�jJj�F�`f�4i/$=��2�.P�Q!�e��E�z�No�Ҏ��Az@#Q��T��Ն��]`s+�8;-n�tum#$-^��m����>�ñ��.-�D�����	A}�HFs�!+�?P���K[�����򁶡���#s�1:X�����*���t�v��8[���!��3W����*^�k�V�h�:N�lw7u���oʎʞ5Y�ª;*��3E���- B���{�rmd���8����ZNl�t����;��Qҕ���d�B��$�b��!"� G���g�4~��2� �o�����\_qP_��[���^����HD0�U� P�1�>E����M�i�<�azT�����������Zo��:��;�!������e+	���[\��'[��R��ѱgg
���RRd�^�=�Dǔ۳S^��d��g̦�yV���������z�I*���8?F�)��c�Ϫ��� z�|߇���?�ump��8�r"!�p�ڊ&�Q!�wA]�{}�lm��:�6w���_Z�!��[>#��bʕ��c��Y��,.v[PQ �< | ����Bx��:_�Eb����S��B���l�jɭ���ҹE_����r3)�y�����]��N^�����ӈ��Ě�<%+��9���p>���������|��q��Mi,';щ������I^�'�^-'9"�	=JB�F�J#g(��d��Jr�mw�q~:�\��[�~u��Dӥ��y�0
R������Q�CsTf�^�(=+;��k^3�(�|5�S��,�^�Xx�};K�j�m]�mr���c5'�\m'A����P!����IE#��zv���=��[����$��������O.�^��Q$��J��^��	�_Z�>����U�)�(en̭��5��ڭE���4/9B���&X�˫�
qj9p���	xqo��At,���ˇ��:)=)��\:*�f�%9a��.֗<��rF��0��h_+J!;\��j!���1�t�����*!:A����!���h{z>���B���K쀱~2��c���wv���s���0^�%J��🜞^�_�u��U�hh���cH�~Wd���[I[Z�jؼ�������J��^��c��R~n\'$̯���!H�P��K]��C��'���Qo�ʁ�wfԬ�k����zRZ��9��_�?:"`�s���~�:GU �uѦ1�,_	H��j�,�����&��[��,�w:����aja��14�/��	�!���l_�^J��q�S�Ǐ���\E�#�F�-כT4ur��8�I��$W8�,�Ȟ��M��;ie��n&�6G��r��e/�/��:�t�T���Q5�5�P;4�sY��9��:��\��{|_s��~�5E��i�C%
�6vv�������R�T�MM��R\<<;p� Xؙ�ZYx�Ύ�ͨ��NB��n���&XBŝ��T*��ݢ�C��,U'��Tԅ�<�>��(t&����B�֢IJ8R4APY�� 6�����N���3�������"_M�-�v�1~�ų�B�{^5lҫUG���7}4�&e#�y�$�%�l�bC��A�I��6R�Oc�0Y1}�#�^�0��6����}>��|�   �YK+jaa!K�G9�i�����X��8O
?l������O����G=���|S����+�y�{��ḙ���T��O�[�kW�b7���<M������o��&��q tP����{4%`��s�W�"��Y��O�z�"�ݙB⿎γ]Z:c�o;�f]맏���!���޶���|�quh��z�[$x{�)��l�
ժ>]L�<��:x0����x����Ύ�[F_���,x�qp2�����Ip���W[~����[5�j�����J��YEv�a7���4%�R=n�F��s��/�#0�^9+[�ޔx����"TT[#�Wv��wGQ�E���K���k��ޱ�wV��.���c�z�~6b��΄体��Gk7��)(�Z!=���lͱU K.ujz:ddD������^�1�#<��-[E_LZN��'�D�n��:�_j	�!�Ǩ�w
����\-��ag����c��w�2��שIdX=��͐ֈ�N��x�T�q{[��u�V��mrPw�*Wj�6R���=F4m�7�q�W�G$�S�r#��Y�Ë��b�6������Ȃe�<>x���ł���'�j��e��ں�+�Z�0�͇H����36l�ʹP�K�����K�iψ�
L��'���ž��n+#�ϑ�%�_�t�3[�c]6~]�����|9�Z�	�+蹝�W�)�Ď��v��/����"���.���ໟ��L��p7IT����ʈ����%Ov��h9��x��p�K\�$8�É~(4��:aE�a�l\i����E���ՏO�;˫&��?1�� t��.f���@�vbUr�(��2)������k�1�c�������v>đj��J�y����]FfF��HxK���ܜ���t�:�P��w~�ӎ�T9F�n0�hUo�^N-I��i�x�b�D�`IO�3��) ^��Ak�x�d.�q5��nU�n�p�,'���H��{��Q���ߧ��1�I��Lnk'�\l,פ�0��q���7mH�|='��x~]�n��pt]A��\���3��m6����a2DvW�Y�dD��%���6����w���My_��6X؁�1����P�=����eh�O(	-�4�w"� p�|���.(��M�I9?r��"��EPG�@��I;�ů��� 87P���U�ڡ����=�c�6G�omaҾ^{]M��a��l+�¥�R-���[�$������nO;IC�7F�Z���]B����+���mwwww	��	�]�����ww�<@p��<�=|�����M�95̜3ջw����)������.�qs�I��\Ґ��w���"��h2�f��D�ӹ����=m.0�M��iæjQ�Y�G:)�q�FP�N3i{Y~S�6�z=�/�<�>_i��&2SA�{zu7�%�Z��]�05c��Wx������Q[˜�gFO.rp���r%lY���OG�ɏlg�{̗Ȱ�Q�}��I�0����|�+ɀ�_�̌�kt�"�Sh*�Bg�̣����2)*�F��L�  2�a�&�x���<�E��	����F
��z�Ϟ
O��<�J��9I�蚴l�@2��$�:���)4?tf�#s��rJ*nm�t_O�z�箿^]jhb�t��L�����~���u$�,�o���1���B������y�K��`u�������������s���jⲍ�����ݟ$eӅ*�Ë����-7|||1��6N��D���u��꺰�m=0��l��!�YOmS1�=��"�_r��p6��?�M�S37�������qހ��ɜKa)����Tbggګ2Ш�ÌW�X}�Abw��g"w�K���ۆ;d�E���o��x��e�M:%t��#�!����igm�����a��
�v���q�G��	r�|<[��lc�->I���C-55����8xF�+��?����Q#M��o��n�.v�5٣E}C8��U�T��8w�m��	2,:�[���}l~p�8z�P9��w(�yH;H`�DzTn���|�0����Bg��?Jb����e�˓X�y�`��85��_�p8l� w*��o�Ý�
'�}%]����I�f_L
� t�'��^J��s9��z�ږW����`�||�|�t�!�<�x���G�}z����Y����_?6'W��	�3z� ���%Y|� };,����Q��n�C߱k���Fc�*y����
ی�<7ڟ�����%>[�O�	��3�\�}�?o@�%$;��r3����>=�)[�}L��iZ�@�Sۆ"�#m�Rw�p���nIy����d�1w��
�t5�}�^��{�x������D@h�(f���;����%BNG���$P��h_�M��v~f�9j�y4�R���n�^�W����dK:|\�J��b)NZ��B�yM��v������2X��/�I,+_�i�n����E������6/��W�l�3����A[!��O)�v�h�s@��\a�>^�9/��(�e�H��u; ����|�5 Tq��E��B����
��J#��G
��z���ٟ�
��
�$O��F�-�*����MDjFw�Tm>�9���&>zƟH�0�w��$5��U�S%�C�� *���&��%�x�Vоb���T�X%W^�mj�k�cN����3W��2V�n�j�e����4�������(�Da�)��>�3�@A�s�^j�ұD��#�@���?���ٙ ���+��j.�L�/"��NcB���3���(b�:���.����Y-%̠rMmo�ꅂVߺ}ֆ�:�}��+��\5H:M�������=k�È���O�U�`��C��=� �Z�ky!��?	Ǩ?�[�����o>�;6겴�����:g�S���Q �� ��O����� ��ԸMm�/2����d�o�7�\��X�FI�.�b�Қ��5���&\�Cx������a��bC��L)��t�Z[I��|𶣕�\Ύ�P��iE>O]��!i�)��Ww��C��؉ �*F�h�?Z�]�ag'��m�V�#�3x�b��,E`歛<�(5���k@)�.�QqL�k_[��ɺ]�!>�)AV�X�k���r�HZEΎa$i|y�V�ى!�"Ob�V�>����mӣ
|�uj{A�Ϸ~"6���N-���m�c�G�����ⅹ9��B��r%z�D�����׏@y�K�(�;�5��Z����vϵ�`���r�AyU;~T!��`�ϑ\��!7���=�(Rk/T�%2�<lP}z�Ap�j��b�H����
��8��3��oM4�e̳�Ą�Uc��p�V������{�5����0�Nj��m9&.E�1��T��kyNk������'�z��#$�n��6�N����-�!F�󚠮iHV����e�,
���5un�y�L���cӝ����EJ�b����kZ<��w�"�˅��k�m]E�:�t�j���1ouF��A��r5MM8�?�$�LHX�5c"� ��M�&���X��Ҡ�|b��<��۟��fP�tx��S]���o���k}��Bh����'3�-������@+헝�e���M� �u%}������\���'c<���O.�x��!f���(�w�� u�}c��G27�IS��Uw��+��=t���A�,������	�W�����G�q�Ӌ�p�c�i0Q�O��]��о�T� ��md�\3���s����(�9m5��>IXd����Y���d�F����S.1o� $��|'�������w�Fi�H;�(��y�����%���������f���*��e&$���fވ�_�� x����Җ(��PNww��v]��s�\'777��,�zk) �	;��i�;�
��Ѡ�%N��J�}�v5�� �GRpxh���4���Y�H�]j����\vдXxt�h�Oe��Vs��q�?AN{k��iq�����+4nS��Y��ڶ�^��Rl�'�Dj
�8���?�X\I_>)����*}��K���}E�_;ֲݟ�N�|�u�w��v����i�Ae�n�,�_[�MY� ��*]���0����F�OvN�Xh͒"G�v#�z}�K����M}�x�:���:\�LޗF��g
��&�v��4ȣxq�p��s7���թ�����6��-�/^����o�d"H�}���0=/�ϊ�����[ ����o��?W$�/��O���qV�51�U��Cp[Gp�ى������A��=QB �غ��> B7����'�U�n=W����??�!�0)�ݸ5@�wY9!x�0l���1:H��l,�H��� �J�hn��~��������cn �O��M�4�3��5b��5�)2~,�	��`{�8��Jk"7��R:V;t�JW���B/�1?Km`Ѣ"�I���]��@R��g�S��۔����GE-�W�L4�z�%���z�����C$�Q��mthk�ed�[<�����4M:���H��7������(W�S������j��T%76J	:��"R��k3>}�e<u;�@C�eGG��3�;�ܖ��0����aa�Ez]A��ᛔܐ�r��%����TW�|
Re4�q���q@pl�e�͊Zs:ކ�u�!l� �N͎��FK�U�KIO�!���>�$R��gȺ�KL�tB��-+���^p-�&Rr��c����b
�[�X۶v?{���Ģ��,S��y�8)�u��	�v$�R�����<m�zs8QB��e�8�ę�p?hN���#!{�������&7%���zE,h�0�W��}�?�����.8��.�5h���3��C�C�ο�������z�ɩ"�k�f�2�!醾!=O���EШ�Q�Q���n?4�|�~գ����Y�r�C�~�]ÎF�{/�' ��.����-x��3���H1���}�_@��E���yqИ��+p�%��!ʏ�ի��}4��ݯ�W��>U ��)��v�o�z>c�U�W㑵��>]94�@��	�b�z���E���F��,��	�	�����I���T�8����`�?���/* �p�7B%�
D|t�&��In����ې��!r����{!!{�!x�4L�z��^�||��*�rz��E<ډ�7�Qz���.:
�<�ZZR"�����̃�O������ϳ�	絭nq֫?k՗>�c`<�M_K�^��'��vXwn_�d@�e筪��ϻ]���[m_ݞ���<�QH��9v�+�vW�����j�p�
@b߄|�A	��n�����f��2����@6����2)"ER�xe���;�j��s�|�Szs�C+��)��M���QZbk���(b&d�r��f�e|_������U4+x	�\X�W��X�"�.v�I��q٢����~�B./a�jp3M\���7�>�,4��teJ^�)��F~�7�5:)�4ut��D�#A��UU���F��!p�Yb����q-_�d^��
�	�p�T���sh?���`��tp1Po脚E���}�R6�SCL��1�J:Kt#O�~�[���E�ɠ�c5��2P����e������,�ාb߹�閭7sQ��!��Il�9b���A���*��GC$Ⲛ��� Bm���.H�P1RsZ0�b��o�J�@�)T{F��|��#��u�	ߣC��`�=�<��گ����6�򕶤D�^*�^y[|l��7>�͸���H���87�1�gd/����E�i�_6y����R�.��b���T�_Bp�4P�#Uf%$�r��aGbU�%!F�UoH�R����W�{K��8VX�VDL("Pn��ku�k�sǷ��Ya��m������BK|�Z���Y뱬(X���bnb�,�{Ǧ��ο�� �d�I)n°>�46�agt)��ށ�N�~�ƫr�Q/wJZ���}��W1�hѥ��EP�2kYfp�o�����^aQt�
<�U�	_�$%0�6�K��O|��Hγ��ư���n7X���I��Ƽ+�'	0�4~3��3K��j_�n2]�����e(��`"�s3�x��O��>�}���FU%�
¼�4�MT�e��䏇���q�9��*i���6����w�p�'3�Ψ1��N �P�g��lK}�F�����;  �K��	b��2���8D�c9��z�d<������?66v^{��U_�PbZ�v(^�*2e9#�h��Cgu=G�4:�x9�A�٧����ʋ�y�6�7Nz��B������q/
OF��>�B�%~�^��<�Y�=�|�~��E=9��r5.�@^Qu��{�Bmb�S{�/����O�&u��R�3s2�E���|k�sk\z޶g�Eav¤�����z[o��N�-�����Bo��y[f�N�L�/N�w�L�1}��;1l����r9�&u �Z������-�NN�C ��r�o�t�s��ح{�~`@�磫���:gKҿ�H�9۽=��i땧-��Ё��WZ?��j��9H�֬�������Y/M
�1>Np97a�^�IZ#�܂��)1��]߅\g<*�NF�i���ѥ���i���		��~2�D�)�|��O#�٥���g_p�!�{�?
xH�*mq���X	���ܯ��ٮ9$��f2vh<�B�x"o�&N�|����]H���Mτ"g�ھY��{t\�j��+݄���^۾{8lz�Ţ�����6���\ֈz��r`橰ߛ��a4���x3���w��f������|7��_x��Hm�Pj5LE�)3֣��bF��buQ���"��jI�t��a��jZ4$�_��L� �&��)@!��V���� jG���D��\W8�I�H�'O��J��P�k��Y��5&EJ5O}��XP>����4����GX�7�4�o3(=�<����&�ʽ��:�P�4/��`l�M�Ai����5��zϿB)�N�yWRKE�2��D���UA����!^�
��,�IL�U�L���AA�))>�:��O ͽj��������'EM��K��y\��z`i�]���jvB��I�H2���h)b���cU6�fI.:|���H�Qfǲ�ᗱ_P\`ɡ�q���J���%�#Ѻ��T�EZ38�����m���В�fu�4Y��;K��U�����<�A�V`5+�Z�Tq�g���-�0����|�3�%��sdddl�	�}��������2�H��� �/�DZ@�RH�_{j+84�vT'h�g�U�{�.��L���"|��O%b��R��x8$>�%��dUN���� _�y�4��i׉^����jk	K#���G���D����x�'����S�QP�G�zoTA>�S����W����Da�96>>�B�38c��J��P	
}��=9<
�P�E@΍�vƢ�w��	����D..[�T6��ZF��M�>Ԛ��30��/y���͸w����|�N�X�?��D���S�)���tݔT�t~�q�,P�_^M�d�q����p��Ɛ7�J�l�J�1�Fl΃���Q�Z�}sV��/��&���;�� ��V�C����A���֛LD�ԏZ^��`�v5�j�A��0��,���J=��>�I|^�]׿�49i #�yA��c�К�!���ԛ���mek29!��FWW��n-������d{�^C�
�M��d��d�L��C����]�[�3!@�������JPPP����D*����Y6�R�"�F-�O�p<�� ���ʽ�~������1��ߏ�@@A~��=�8��5��ɽH�w%�A���u�h�͝�s��8��Li+]گ��v\��Z:0���4t\9�e��y�;�!f"��n��Ҧ��M]co�΁�Qf�� IEe��^�%:���1���=v���P2�z���sR��,k�S���oi �7#�"5���yuS�����qk�h���l���b�2@Ĵ�/C=��͠�V�v%i�6�H�cه�Ͳ�� ��T|:I8��Ii�9�B^�ϲ W�����������#���1�s>����q�c���(�m�6��~����|�DlԈ��"��jw5f�ez/���;o�#K��ϊ�P��}<,''Ǆf��@�9���>8�6�儞�M�����9*﹗3�����������R��W��7�#���1���q`(�]��JB�_)�&�ƆtlJƒ�aLa�BC�\��$Zs#�s���9�ⵯ�3�Eޢq4Y�)�³6DTGe?`���p��ww+�����7Q�fЎ׻��1�9��%U%�1�ͰO����.$�Ќ�6n��~��37�9���t�w3�3�|���u�{��g���9�0����� ��i��>��i�D1DS�9n�!vc�:D|�gmm8���4�@�&Ad���dH��V���u�w�Avw�6���+	��*�Oϝv�ϞfV$�a�ӬT*;���w��3UD/0�Ư�
������-���a�������ׅ�i�O���g}B��G�DE�ϙ�t���u�)Ն���>���uKិ�	����ذ!�!���7�?M9��#����Ĭz��eк+���[��Zj�>f�\�9q>"�"|�`��UB��zOլ�#>�|�STDqh��������%��L
'ӛ�� /ݙQ`��������~?�*�Sd �]��KU�5�G���:�k�U�������?��!Z�a���Q��2/K�7����+(n��h!:�M��Ȱ�n����S:�_��Ϝ�'V������@����#�q��RQ���yО8�uC�NN�Di"O�K���O�:�q��ȟ��(����ơT���,����Դ�=]r�/(AHfFE<�����*3ȋ��t�<�la�;���XX��LL0x�������*���;!�}S�`v�@ Z v�U�q.����T?JL�]5|�d��c0,��PF��<#���� vX��w�\���=_�ؾ��ܒ5�ǳ;���v����"4��9@�	Qީ]��mJ_w��%�o�)�v���Dk� �DUB�	W����.ZY�0.������Ed����~ ����5Ʋ�e+�/V*�҅�>��2��Χ��v"u����8:x\����(@|u�����X��C:q����J;E�Ó�˱�]H��H�/��U�Ս<o�D���Y�t����t+��)Z{{;�W�do����ӞI2���7 ��כ���SnaM+h�wa{a��d+x`M�>M/��=`��|)�ʯ�1�%K����d�����g�b��ז
����]U�{PZ>?0-c|@.�M�%a\zVo���x�v��#��� �<�=�'�|�xUv����%�t)�[�Xֳ�~�'�I(����.h�64V+�XN�b̋zˈ�)���@!`��ŗA�x�:����`�;����贪���=�{���;vΒ�Z4�e���Lpp0drrr��<�N�{P ̎��zS�������Vq���PԿ�ݨ9B|���k��wg��3�TN�
z�-� ��7M[�+�����]��5f=60w�`�\6�B���K��y���	����w)%mIky���<j_ O��i�d�E��qU��@f��/��c��)����J����^$
���s��Zc����pq��Q��� �[�N�-|m
��x�$����<<vD_wE�nU�66��Ӕ($B��� #[)�뵬�VFCc��hZ��\��I�yV��>���b�Bs�ej����<9�P{|WP���B�͓�ǉq��9p9�5������\@O4��^�(�� <g k8�˧`�i���j'����)o?��(RM��f��$:����㛗��p�C�W]Ԯxk�G�n�����T���Zt�l���>�#]V_�hFae``>����kyz�{��v/���[��U��5���#�Ѣ�ȡwvv|�?](�����Ϳ���~gboo�ߛ�h���+_V^.�.b�����΋Ȅ)�0��|��X�~�p<-�Q���#پ�d�xr}E{P���H�ɱWH�6��Wi����'�$�Z�({#�/����!1�F���_���A�5��'>�!Htc'S�o�J8���H�)/���!�Tɸ	I���:�
z��ja��4����=};��aז�^~��V�ᗃ꒎�u�}���(L����Is4�D�&3\��%�����zZ���ӟ?�^�[���u��8�Pz�y<>2[4�8'd���c��`�a>]x{{{e��WG��!�9sF�}n�}ؕ1�Rh���BUW:"��X��A��d=�3k�� tLZ�${�8<�������F�E�)XhB&�'3�q��H�a�[�
M�k|y���54����z�������>�yv( %�؝cys���z�����C�����0N��sT��:���'��Y��*��GrYQ�_1��'Y���-h�R�����`���.j,$����I�U�lD/���M�!���L�'F��o��2B�u���T���j����5D�(ihH
HWNc��,�@�i=�tH�r'v�!�s�5�%�Y�f3Д���f��/>yj�&�8}���}��f���A�Ű�bئ蒨���K�sy�pB�3:���?�c�9]B�S ɝW6Dյ�:�G8��U�k��B#��>k`D������r't3x���c�������9��.�G~�Z͙����ɟ��^0��l��?B7\����/Y����s/�Ϋ���yd����:�.��10��Zn��ۓ8���F�3���|Dݟʍ�����S�u���p`;إzީV������	�Ԝ��w*�t��:*M�ƀ0�>��#�+��-@n�ED)�郵��v�9gU=ږD]y	�]Hl����g2�N��N,�QB���E��;�]��=���dȃ�,񙲑���Rj.PpF��5cr_N�����r|�����׶	�b�ֿ��٧��!/�^�Y��n���â>T�`pbbb�n>Eh����ˡ��(�O	�i�='�?Q`��D�2��ǑE��ڧT'7Pҫ&�h@�/0�PZk�<)�ӎ#7Ð��s�b�(���&"���� �6��'3�~_���U�,��h�f�!����8o��`!墁Y��H���X�Gd3o�eA�Tpq\���f=�j"�j	���4B�����{8nr1�4�.�����#��V<��s�9]����O_w�v�](�S�[���\����P�x��f��w�VW ���� Vw��}�^a����DJRF�n�*�0Bz'p���s��}�{#���)W���S���>p(�����;�k�%�<���q�œ�kz�!�^�8j��6L��*�����Q�W힮��<�R忷�K�Ka���^>����G4��lAϝ��FC�S�� MDFA�sh ��?�ぁc�l�����]g�$�����'���M���\�:� �1��������$��O/º׺�[H�]U��q�5�W��V�؋�,�tO9ִ�c28��m~2Q�"hHl���D��r��	/��Ps�[6E�c�����f�~��@�5i�u~{�7;���s�o�w�A���v�Ǎ��3n���Y7�>��MM�fQbCet���K�1EB ;��([}ٞQ��<��턉���)))��J�0�<۽��3�I~~yYs�.2��*f��_m);t�etl;D뉮�U�r�^�ȺsV׃�I�M{�`��0�k�t��ž7�'@�߯�ds�y�T$FR��*J¿�L$����E��%�B�N�1��_��?���=9������R�ԑ|�b������ѐ�D5��M��nGjU������������u��T1[B�eڟz�LDQ�ז��z��]ҡ�1�Ϋ�x�tʞ��_�����ڙ��]�v	�V�P|)N�H��<��p��#q|�d��2����t�gl}f*�j��X��������gE�%��Feuu�a�0q��W �aX��Qs�>c�f��p��:(7��-�w��59����JIO�a�"��^B����y55�>| ����S�?�ճ�V��Ċ�z�\��/�b�T?!�rN^E�H�Տ�a:I� �i�40�@~�Xŕ�d���Q�hs$�vb��Řl�e����)�w�y�Vg����K+�HZZ�K��j���3�X�SѨ���1��j<�(�u��2��� `������<����4�#FM��)h�T�x�g<�����!���)�F��!��z��Ly��QU%+M���,py�o��,3mS8��I��JU�?=�4	�8��"zLZB��W�:x�������q����^����i������)G����g�I�55!A�5�8�%S�+*T4���p�u
��-�UPPf�b��E�:<��(��jf�$�/���a��&�Kq3�����^��Z���6������� �u3�7���"����$lmTg{�OG���e��Z�y2�y�_��Q�q�qwx��$JB����n�+8�xՍb)�}�gT�F��k�>:w����Z���������w��ON�>�!�k����%�A4�=�����Ynn���~"df����(�#���؍Fa$o&V�3�	F�َ[��9���!:
��yo��y��0���|g�3���u�*�N�a��>Ƽ9/k����sS������3�ǁ�F���Q<h�.�=�nOX����y���;�'�{�	�u�]D�K�\$
�e�K��Z�*�z��j7! 5l�n2��ď��^;>�i���21_� �j�^ ��VS:7A^��r�3�7%�?}[�F8\Yʺ�TK��;f����a���%��5X�C)��{��_p���)�HG`��S�ۖ3�sE��[�䷴I��������Xtn���"�s<�҆��(��|=Q�!X�ń��q�l�����5C��tn�b,ŞE�=:�]��:2e�Qlh$�'?~^�-O�CeK}E9l�z2�~<�j�z#�jopF4fcbddd�^�J�_@>>���=*?Ñ��tzG�ab`�:;C�
$�2Q��4B??�o3��`�����4��E/8Y;ڠx~Qp�~{�#][�s��-v �Ƙ0F&��6;&k�b`L# �||�F���U�t#Q����ǧw��:{�y���-KjXtʂm�liv|�c�P��&��Ev��	��&N�ay�o8��*n`��.��#5ޠHxpn�I{���`L�Cx�����8��@�/v�Ah<��i
F��\�|,`��S~:l�T��%Pr�*&�:P�2����ôQ���j����[R�	$%���$͓+Nc\I_n��me���xC"��w��)����,���h�Ca����QW���8bU0jfY?�!:D��������=������9E:ં�H=5U�R3�>�����`�ʼ�N=�dO(ñ	��q �RkW9.�4]������r�����f�����e@W՚հ�i&�nEݣ����{��ڌ�2읙��������^v�)�9��n��y�h��Q_�-(��fT�5�Iho#0��x�'�n�إʦD��L�:�Xr��GHt��c�U����Z>V�~�ན�<�]E�K�r��pi����
e$�4đ^��K���js���>*�Wڕ�B���w�
��I8o��)0*���1�t�eX��2�$���/4�t)�K�_q߃5sJ>���.���������jXW�?�>�D�ؠ3t�(�"��uC,!r맰��
���UH��,F�g��\�R �Bk?}�ܓ����|�N�������_��T��o�5ۢ�(5�'"�t��U�[if�^B-|O��~�?�ǊzW��AtX�j��:��:��-������8��׵" j�(���Y?��鯇�,H�g��� -�����˞�j��Q�^M������P9����:��3��vG��
��*��r�ݦ�z�D��;V�.�ipl�R�zD��΅�7�tD�w!GH,p�eT��/v@}ϸ�O�nk�L�&��?�k�S?7�}<Ԩ�Y�XdN����l��-:�����<̾�"��G��%t�;r�̇�fp�V�oK*�b�;.�7��Rih�Ǧy*����_j-�U�@,��H5K4h�3&�!V����P�ˀ��^��"C�Jo6xć����y��Ҿ�~2mr��s�^��r?0OR�-�ܤ��;��9b���Ft�$�\��F��@L���J�M�JC?A��q/�7�7���6�ժ˥j�ء������*����M���	��_9-�P���-/j��v��Ư�����Z���<s�kD(�@��p�:}�5�sE5���\"z�V�B��éu~�Y1dTIj���Nv�v}�f�</�nO'8H��.�g�}�S�6_�L�Q�I���c��O��;��=�:k��Hd���x�yu7��;LKe���@�TӍ�۲2�`�4AZ����~�,�;=��Ǹ�����%�	�x:BZ[�.�Yp�Y�#c'[�L�/AJ��H�g!%{�޴���x���	�ZF��������ŧ�2~	|ݗ;�Wq���'����&���)�=��&숃˺���r�������kד�����N�;�<�]&]��kؕ�������j0Mf�Ө����o�+��_7"�6ɪ��>PxN)����z���=�W�r��<�:�:�N,-��l�V����.a����ŇCR֭]�Z�v+�2P<�SGYƕT�����d	�#�;<s��nu��/��(i,TA��P_	��y�jV�`9(�9w�|nC��7�깂:<�y�����F_zot����(�s�a�4iJ9�{�C���fe����G���;��W �=s��o��pD��{q7��oGz��>\Xv�zY���i6#��6�}M��7C=�X�z�i�}	�L��C�,�.R�@��I�"~Ґٰ�s��mU����:zh�������Y�Ы�Ԟa��fD��$��r����}�*�~SQ�Ϊ#� ����9�(w��GU�F�L���9��'N�f������߽�����[�ڝ5�CPX;`N5�b�㢻u�ek� �*��;��%�����j+��z�k  �����/M�a6���U84.��g��/�{=�	|�6yF#w��2z\�ş~�T��R'��I���Pz"�AH$�1�H��/�8,ںF( �����E�O�)�^�6�U�	�;��k(_�M�3$J|e���d�[NVd�-|]k����u5Q����s�)���P��;uD��Uj��5��v?���n����ا��[�RS�7|A	��1k{Cd�ޓD���s*4L|خ��q�؍2�cC�V�y:��6��+����k>�b�G��)�hh$(��WC/�����Y{�,���)ښ�q��t@Xkf:�i�P]{��o{�*:�|@�?��>��:h�*�v��l�h����cGZ��տ 3�'�,���F�Q�ۼ�����x^�p���nE�8���c�`m���Y������X��C{�ř����[�&��T�����틳X#�O"��%3��+*X�㵩�ڿoۏ~����5b�`D�U�������<:���[�x�^�{R��.�����ѹ; p�o��5�����WO�����Yv1f�_��,Hx���V�f��������x�tL���2-lX>x�W\�^�M$\1���>&��J�L_l��&�f�'1$������=�P��0��~)]a$.c}(����ȻmV.o������v��#J�!����:��M�o�o���||	f5n�B7%����i��}Y������iv�MD�7�O�V,�Q�4��mڢ���@6��wֈ$D��&Sjm���1������`9�S��l���1�g�'���4�$� ���wK�y[C�~�o�`[دܱ�~�?��D��y���j*vԜ�e�t��8'��s���J5~��޲=v\���~uI�K֊�O]@����u���G��$;�x���_�!Z{B|�������TPK�$����΃�y��d�i�:��R�O�xlwzL��S���~b8��]5���2P5��b|���Y��lX�ST_K>A�Ɂ�+�
]��f�
��FdK`u��|
f��hg�B����l���E^_7�[�\��xz�H���:���^j4��k���s�g~f`N��Z�^���´��r�G��JU뾢��D:S��;{�4�]�B� �3���p�[Y��&�j۔Q����O�VyT�yt�e�x�x�jl�3F��{������ߥ�s5ǟs��	���P{�ޢE�c��9Mf��z����f���/�[+p��A��Szaw?��A�pa���n�ƶ>���i�V\����o'�k�E�W�&��e����)N(�d�Q�rL�Gk_5s�iI�=}�載`�`�E,�N�%��]tw��矶��Z��_&8���<g��[^@5�I���O~�t�6O��찶�\��=}���7����uq��o߷t�B5�z% 8?_Rk�}��)�c�ZG�1�����`=̇G�\�=6-����"�?���[��ݗ�h'�/�M�_B�h�N_�����A���Uu�T����"
y[Ջv�iI�w�b��g�堙���g>Oo��kM>ʇ(t�����t9^�"�k�52�o�y��?`
�?�q��K�)��S������.&<��0]�KB��L�Q�ve�Y�����ԸC(5�g��Y-fTpN�@79������xg؉��%V������6�=���h)XǢ�=��*P�}�ir}�$b� ��e�\�3a�ץoG�/�R���/�'=����9��ɓ1l��N�X���7SO]��j�p�6�j%����2�T��W�?��G����I������bF�nzH�';�!Lh�i��:m{�D��M�,my=!*y��x"�v�/�:T���,�;����4���YҞ���p6�mo���o�z��[+��˱�&n^����M;���/$0��B�b�C'[}�.��Q�2���πS��j#oB8���N��~�S�p��xǒ"K�p�M����XjD�����6̑[{�Q,����M�����<3�\���@|����������N��*\�(������R��gC(�J�3�d9�T�~�U2�l��/D�?�5w �GS��{x���69��۲Vdol��d�qS��P��RCX����HW�o8�7�=*	����W�>���b$*wpr�}_u���QE2-�Y�z*f���8V�Q�&�f?���OǗ���d��4�Dsz�%Ζ}�Af�_/�#�S����R=���+���F&��1fx�YДe��tF�FĂ�/����:�ܤ�@=υh�FF��=μ��6O�r��}�Z<D8�S���5'Th�3-��	�tǾ@�d����LpWD��ՙ	��)k�H1�	m{��cWr�u_{���N<��+6�l��xw�[g%Y�k.�VR��V��&|�<d�Ώ�U������D-*1�<�,#�7�t4�y0�a���ʲN|u�lI5��lL��~����ͭO]	���S��>��V��=E��m�Z��}68Ǭ6L�}�����a-_$F�3��W�Z�g� ����+-�T�$R&xH~_�$�@h�!iQ�e�Z6v3GJ'좊���WҢ��m���{����-ܠ����{�*��Yˮ�:�)����Ӊ�?��K���芡��ۭ�,����� zy.�@� ��Gs�+C�b����[�hf�x=qZ��^]�'�/�$����}Z�_b=
�I�ژ,}{>`���TT�cnКɃʿ�|n������L�R'�P{��o�]_+Z�AQ��7�ny��s���t�Ã;���!�wwwww����݃�&�������'�+����a�T�޽W����>5��b7���Z?g�켯>m}�$;l��G��qo�O4;�E#>��r[>��w_�h��b"�Q�C [��[ٻQ�D��⯖W%��u�n�h��	�O���G���D�Y��R{ �,~p��۲���z�Ğ�W,]��=w}����{�f�W�]Ix��6���U[��5���gN�!6=���D���\��� ��O�I�@ű6y #��n������60P>�wt�F	�!�j裂(�P��;�D���ި�������\Kџn��,��u.]�q�f=���=7�fQ8@D��A#������t�}rq�U"�	��1�/��a7����l'�3�_�ZGn{y؟?H�}o���u���@�/B$<�r�m$��½���Ih%ڳq����%�ɢK�43�m�y ��+����m�v�/��X�Kc LS�=���hIG>Ǹ �j���>�Vs�����-[�SJ}4f���w��ݬ�00�&����ȑcH8}���B���&M�����&D�9q� �~�Ȣo*j�Y��df׷�K������zv�:��]יh��!�z%���)��v������p4��<.��YD@E�(}j��y�ג3��s� ��d0]�q��BF�tq�XSe�s���1a��J~c�'�]l}�=�jh�(�n��j� ��c ����$���,Z> r�Y����m�?�l��3���$ad�;�aQ�w *�e�>��Z�� ��~R���1|dr�}�)onx�?��^��Ȼ�T}߽��+]���'Տ۱�b��s����!���m��(���pZ�u�e�H�9�W[�F�P�������JB���N�3����7"�I��6Cn4y��n�G�8�|�y��|q�a�.�y˸'^��Ԏ��{��о�VB�M�hb�`��}2�6SU�u�1 l4��h��%�{�>���2m�Hc�l��F����F9+���̲����d 	~�̫�3�"ȝ08/�Z	���ʱ��W�OZ!.W������W�Y��I�f���H���@A��T��#iz�k�t$�����eVPh�y��\ �%l��h$����?V����	�j�B%4���z>�U2�M��9��XI��i��m\�x�:����Ā0��m�hv����⺦��O� �]&��~=Y��f7��X,�:s(��&�i���؜��#��:��"�*ǫ�OK�>�O�͸����ZI���>J�݂@5�x�6��J�^J�\�K"�1�e�M�
c0_�j3�^����V_�D�	S�7J�1R��ń�]&D�q��ڥ��jrw,��t��|�r�������sPҎ,(�u&�	�c�DM�j{Q`���wt��a]i����j��[Eؕ��+QVÎ�Lr$U�~Qm$΁�V��U %"3#��o��Q$.�Ly��bƠ$@��2��l(!��a���;�c;fN���}��'��LN�ciwÁ�������@G��~�jO�7ƚʬ��P�>.�_�r�j؈yz5,�͟Vw����$�{�T����Yߖ���,#"�l��m��2��o!.�ӌ��G��,rOW�2+�P���jԦ#�V:��j�zЮ�R��}��&�(k���k���\�s����5��'_i��Y7�mI�R\/9�F��>V���>�P̿����x5��	0�	(�{w�$	��Go=��*O�y��>j$	`9�"M��̼p��D�ˋ Q�Or��QR&���3�â~�p�d�V� 0:�Bo�[�h
>4{$@'�F����|:�>:V8K��{n�׆:g>qz�By`�>�^a٧+�q]����[�G�GM�IR}��G]8Tl�����ߤh(�Q���U�"a�1�F���PB�p�e:+q�j؅J�����Ћ++G�
Nf�Y�5*�3<&��p_tɍ���U�*��mMvS��k�>��I��u}p�
n�Vt���Aa���]&Lц�GC�:%d�Y��;��˷�������{w�z�
��O\ywJ�o��3f�������#���#���pj�Kt>��f��\�P�X�L���zҥj���YY��1�,��L�4f�cG�͞��!�7#�m���& �`?)�!ڜ�1?v[�,�Y�Z�
�<�ƴ�y�:t�7��/8k���M���p���**(��CF/�q}���O�)ID�M/���Ǜs��A�&���Jo#$�]��($	��ݻY9��$���n դ�IE�sC�O��q��q糶�49������� ���9�?0���x���������z�N� C�Y�p�����I��~{wYY���r̰qд�-�K���F�ۥ����ok�߸�n���ͬE��k� b܇�%!��OIR�ifb�]� M��F��c�
�T�fs�$@�iXM��7T<>Hy�2�d"B�.T�~���;�:[:�������3��$���H�Vpp�]H���=%wOFR 0ٰ�
�u�yv7��j�#J��Ng��I�st�륈De��ԝ�L��X$5���������� 9 \�X�
�Y��0���})�++D��/l��֪&̡L�Ύ����7� �cD	;m�ޖ	w]��)��%׍b׹ݣׇk��
�\��e�� �@�Rw#33Jq��Y6vv��Y.;Εxq
J�Z@A�p>�|��g��"C
���#@�<<��-2@�k��y��{�NdEx������=2[��>�"���U���\�;g=��^9p�.Vn^v|��U�*��v̅��SU�)E�$.j��g,Dl_�|������(Oxb?fL/�s.�����jI��=�����S����9v��1�~C I��uWǷ�g�ӎxZ�����fe %�����`Aj�s@��8���&��#�ƪ�pnC���tQۀ@b@�'hȓz����_�Rc�����\��6��~�C��6�7jY����\�0Km��^���o�FG�'@`��~E>2�U������n����?�;�f%,l���OU����_����T��~2����'�AG���Kf+ʣ�ҋ܆�cS�����I��%����j�f���������1]4d�N��+q
����&n0�ҙϹ|sӃ�̹�tQ��V��W��>6\���zCy7?2�rn V��?B�ў���aь��E&͗q��]ӫ:�@��5?	�I�L���>r���\se����q����@E(�`Xf�J" yQ��j $u�}_�t����QϏ���ŝ*}X�H��e������&z�eii|2ev+`zj�ב6���j�+�έ��vB�iw�&��s�ᣀ�H����'�q��Y�A��}�YXu�Q�v�;A�x�Y�����1�f�+\ ���	;,ܞ#��+�˶�}����6�
1�t��Z����M%�d�ڷ1:���2�2�X�W�#k �UO�rjk�*.�fJO�
Ñ7W"� ]�0�k-�= P�?� � �O�=��O���cwY��6��̗���R��V�Kx�h�[=5�Ѽ ���>�d_�+�Y����Mӄ~sC����<�:MیnÅ�$��';U�����y#6$]t�8��4kP�R-j��g����PWCS�����;�����l�<V��vsJ���b�G�)��h
?����MU�)r��P~92(7��xbOԓ�7���(0��2H�|$�Җ�i~�����^!e����	566����O�~fH)P��O������V��6�����@�f����Q]�ME�ܑ��η��L�A�<�Rp�Rm�Q�@�
LQW=I�T��|��y�n�����yk)v�i.&�s 󱷋���:�������tA3��8�>!*�Ĩf��p[�J��N�Ξ�͞6���t�3e��#ƚ�T�I��m�ًf�v~��C���w=���Ҧ��ug�C-)݄Hv?SN:_�-�s�Ud����~O��ܞPp��z]�(v��Ŗ��ǳ�s*��<��5����4iVm�5���'�����C@t�JA�Ƿ�-����NK�7׭���Y���eS,�@����}��$3@�p�_Y�>����5�����5ɢ)L��\�d��3ڣ��� ��ᷴ;���0 r���,te�N�8�}?���5�0�5�2��} �=J��y=�y�b��vM놻ǡ*e��#����M���J�40�	�9�4�žzt�A(��!���={t'�qfw��{��M�
�-��_m#D<?�1��MpTE��44�~�`�R^p��I�w�\dB~ȝ=�Wý^���c���!��+�VQ&���bv�1�����#b�,^����t?�ǆ�&�a���K�WE&&h�l5����U  ���q 9U_�M�`
�ؚӑ��'�]L�'aU��f��\�����*�'�2\`^`$�w��>:E4u:��-�L$�F�--S�6���z��~���!�A��=����)xʴn�ɕz�����0P��I��~��˥\�n�K�4���`� ��k��e"z���{���'��͆zW�A�]�N��U%�O�2�Z�Q��(b8���In17{�1�G���_ T�yB�8o�L��s�g�!m�B�����Hq�E�T�_Ru��t{!o^����ե�G)Ä����BA]+A�Ct�M2pE#FX����(~�˴���s�bQ�-���׀� �
�����?280[;�c�G������
�h(��p��D�o��2���U��T���T��)�e�P��\iݹ�S�`����QN�"�Ӕ� y�ڇq��җ��ZDT� �'���őۏ'��� �'�L��^XȄ��cFQJ���5s����R=����	-��~@]56��.���bd&��(fE���Y�@��F�@ ���UƯ�#�.j@��
&4���w�߽c;��˓��'-c�w�a`BDb,:a�?�3���y�W������+�*�'EJA�6dEQVW�a�Y�(�aN��j��*�~d2�t�h�R*ּFV�W~q~�HOvx�I7��'v��i�0I��`�U��A��7ɿKY ��q��~'2E ���;�EM{3��������&{�.sƮ�e(��@xT��@�C������;��4���SI%WP���F]zZ�5L�_k+z��N%~�3A��[�8�{M܂�x�k �¯2RpJ���X}���XW�d���e|+�W�����_w�I���/�=B����˩�C�\�*���ږ���by3�œz 1l�@�4�@%2Z�a{�|�gU�}]�ݷ��$D�2DD�;,�D&E%�^m��wD:��u��m�����&U� �'K7�����23�z}5�h�(���^)]��[��'`����{����m����9a�j�՞�����/���/��u��-ϖ�lQ`��|���8��9�x��BL�P�4�.�x� ކQF�JN�5�U�<%죙U����]�"�� iN��C�5�n�u,ځ����.eD�˩���y�F[����OV���TM˄ԎO��]�7{k��T������Z��I�4{�!]�7�k[s�M��0Nd��/|>�k�G��1Fs�Q{�&\	'�
����T���&�_����:y���:�9���n[��t���5J��a��dS�XǼzA��{��Q���!!_��?����U/�����!���ҵ�U��Ϯ�LmQ�ĝ港�/�T�ZoX3�h���M�
�(��V5g*�iw+��Ř$G����P��F���`t>�`��;����A�奄�����t�x5</Κ��KX�z���F;|9+���*���f��	k�e��W�2�Y�ʺ>�Q��x��.+ף�)
D���Sz�����fP]�=O���ּ�;��1-�;^/t����W��<�w�=`"J�4��r������!BMA��B���������J�$w�	�?�iW|��a�kj�x�j�EX����9>�������7�i^G3��i]�0Epeg�q��V���p���փ��%/�:[eg�<��;�o�7�1�E����_e1n/��5S�V���*1���ԛJϹSB_<喚2�S�"��>�!؂8�9U:Ci(~DEZ��V���k����W�,q�R$��u����62t?����Y,�����]ɐ�e��u1UW0�m4�QR��������k満�/R���	�}H�H�������߀�i��Q�d�0��F�"
�L��a'b1 ߸�|�C�I76Ҳ��N\\շh 0����qft��O�~�VOar��Qj((xtt�Y�=���H�Ï(���0Y�D##�9?:��!�w��������kr�Y��
�������HD����u���p������~XcM��ˆ�]Ƣ��5��k����v"��5uT{��Q��_4č��:CŁ�I^\3��b�UA\�W���0f_M>y�_�c���?�~�byRc���Z���_�m0 ��c�hR�~f-w_[���m�βC ���f����w��z����Dx�4��9�¾j�,�h���a��`���pH(��"8i��A"ZW�*��&7��|��Q�D����L�23o�D��M��D=�xFˎ`��N��Hw��8��<�B*�olɔ�PT�l��Zs/�0�-�-�}�+6�-17�ˁ� O5	H1��B޸�!Vm�+�]B_Íᱟ[����o�Y�5��o<@�X��}@s?r�ˢZ[3L�#y�hzV6��.�`�c�NY�#)Vp?y�豂΍L�K��8%:��S�\H�l^IЖ�(��Iu�6�f����5�`d�JY=��P?-��Y�ym\��R���+\�O|����x�x���"����p������o3la"P�����/TQƽHIΣd�W�ح�Ș�1U���Cd�e��� ���`�.x�B�U_�b�9��Z{����y��z�z�.�d����Y��@�?G
���u|�VO�CUGЦ$�*Y���}{m�����[�ǂ�;�5$Hm��ڢ d�}�>D1�,`6���3� ��(? ,�h�hvˢ���F�e]�aH�\�������|�,���
maaS��<y�IU.��������0v5_���ݧ�d	q�9v$R|drqӒ�x:A�� Y���1��(u�R���.S�:��Ҿ���4W�Y���Cl�EVF
�U��^�,;�a�����"e���~r�D�X�E�0x��1Fb��xvA�	�֭�&�R�Cʫ�I��ԏ��C���h(J�<4?�O���,�t�90	�,�3n�SVY	�f�����v� ��͏+)��DB��:�0x�s����хQ1t+�V�YVl.�4fO������RQe/�w@��2��@�ؠg���s�s��|Q��y�PɊ�w^9:�ve��´�2z��2����y�߁���9l�0�K؞��
˜�,���ۈRW6���:R!Rd�qqj��IX1x�ߧL��PN8#o��AV3����4#+}��`�iW������ks��z��L�f��PR�A�6���a��zl�1iۡ�[9NଔQ�?�
6�0cL���y+��I�jd<=xTgt�	�XS)�����nI�Ľͻ���(�P�X��DF&�?���b&A\=���S����}��4��s6ZA@Cq�����S��~�ȧ����}�y匑�"K���䁫�P�Y+�%y��gsU�,y��'W���	^���+]�A�s+�(;@h[��5�]��-����[.����
����t5��a(CL�^'��	kL-�u��$h��#��j��g���:{�p��h��?�ׅ��P����kIL#M1�Ч���g��[MG�f�:���3�����]���6�<��E2
v�R@�;�N�4��~�WM9��PK�qG$�u���0@�`3Y.%7����zt�yd���-'n����4bO��A�Gԝ���*pG]�tD�a
P8:�@����ɤ�mg��@)U��	�^�ՉJ.җb3ԟp���5����[q�6G.�6�&����ܔ���Mn��������M�dV�y/�E�b�/t9�$W��Fz� �+�=�I��v����H/����94�TC�}���i������{��G���6�{`�|��W�	헠����!/"i�c�>�*Z*�w�%Vk�
q���d�L��{p�n��`Q�C���4��dɠ�Q#�{�s]0YA�7�)!na���«>r��bG�KX�.E�~�1�+ �O����͟j��=&�j�9W��D�|7��Ф(�����s/t�
NA�9�S���)��>�[�lu��o���ڍ�bo�wV�?o�/�{�U�����z�.��>̮{���5E��n���"7Ҧ��r�#�#Kj���韖���P��u�˥�H�v/_���uh����m���t�`hP)�#�]4�z����{<�����8���V�}�����p��4��c)5���HfQ+r(!�J��</��O��?��_��;��
퐌��w��J����i��.��H�X.z�<���U͆���y�����6	��m�K��.��NGc�%=��u������ �t�%7A��ZÍ{6�Q
z6N�`����@�J �E}�L���jӛ���,�㬛if�I�T��Z]tb���v���×��ڶM��9����=��{2$�����
)��|L	�_x�8�ѷ[9k���Ev�M2�h
��-�5����Z��KpyE���t��C�c]��}��� �A��/�>\�����C*S�ʯ����)�;p�~m�A8u桝�6£��W�Ȳ������T�t);z�,+��O���������SC���iנ��JE�l�Q��9޶8��{�wͯ~]tf[�e���f	1�^�)�z��'�Vm�
=@^��g�P��6���^��c�:v���kt�~$7�(yE!�$�4& ������K��(����ӳ1wo�C�}�j�'����!F��6s'/���FًJ����_��	��#���7�E| p���kpr�ә�!<��I�������8��R�v�b/��N��p��	g��9ݔ��BW��B�-��jQUɡ^K���ij��#��ֳ�掠�i�P'��?MmE�ɬz.H���{
&M!V�Ԁ�
�ޤJ1�Ox��y]윪��o܃*�q~hu���G���h�_��s2��I(G�~]p���l95g�ѷ~�f�Ao���d�}�����t��Ty�d=i'��
D�����~�Ot���m�5�3C�0~�Ӡ	����E_��q���������J(@X���C��Q��������э�RL�{�pR�?�m����z�	F�l�<g��Y�:b��z�,��z��ϟIٻ����W�l
RfC'N��n��l�O�|q=���9�'�_(���x�E�^��=�}����)M�&�>��V����pc�}$����]�,k�O�f	��PHEz^��k�%|*����	ȗ>=:��4y��9m3$��+P�tH��0��F73ڕvB��r�nZ�Z�?A�R�۞��~-ׇ�����hQ���/D���F������c �4����A���a��*"m����,���r��3~K��t��IZ�.�^�5�d�r�y�U<�cx�-!�����³���/��ll���[�;ރ+�����/���h������/��+S��u��8���|��vNS�����e�K\	^��]Dq+�m�A-�3�1�8��H�hd�����'�cRIW��w��&�������Kb?�^M�5mO_�?Ś��'������I۪�������<��惋�J�
����^�J�q�[�Ŵr��B��[al�r��Wv���ۧ(sי)��?~��M�#�U��ik�*W��_^+U� b�F�#`�n�s,Oy�ӽ�����r�K�"ZAʼ��9(z��� �!}TQһ�K��n��E��e�@�y:W�������~��{v����n�����Xyϻ�3�� f�.�um'��ٿw�����7���Q���UZ��߰�������b���c�#qt�
�~�&�u�&�4b%���u}ǣ��:��s4���Q���ٮ� �1y�+�s���[�<��Y�Y)�Zc����*�᠙��� �:z��N�;��Ңc��ID��Ƿ��7Iy܎h�7�~�7GT�B�q��D����z|)��<_��O~{|٘�!e޽��KB��9�*�_�'���.�|�d�NԺe��0Ns51���S׹���ϫar��
�T��h
��h�l�i���y��4q�8w
^6��o+#����w����V}Z�	k���v���Z4m#���+=e�������̪#�#���/��|}ص�4�x<�G��
T$|f�s�z�2M	���t�����%�����Qҧ�A���MQmJ֣E~jаF,�;��nq?H��K�f��#k���.��E�G�p��ǿS̢�}��4�=�%��9�'�sEm7&�n�MP)���M�nF��p )/�(~h�k��*����FP�-h��B^D�!��ɧ�k���� e���l�A٩�7B���a�N��_�Ub�f��l� ��Oo�\��v>*��h��.��>?"�܄�b��y[�p�����Q|�(_��7����3�=�?�iy��zo`�i�Ik��:1��h���Db��G���8�_��nΐ%���q���������p����:� S����L�ó��$�?����hkϻ�x�󬭷KG /���U�M�L��q�8j��EHv������k%��X�>N��@[L�fRB�J�K"8��qM�*Mx�����mܫ1i�a#�i���[T҃��;z�o��j!)K���1��f��;���U��t�>	�Ed!�i�U�����VR���aV�$2�@8��+}#]u�-]n�����Y��!O�G�)o�����v���p���&o��[�a?ҭ�q�1����9���N�5ѵ��C��6�Y>`��~-�[Qn En�O�[&��I�!���*���&f��?k";��Os�Wr�x�/���DL��7uC�!�2�yLa���pNU���E0ϛ��T�޿�*��>��-x�`\�}������qN�x��	,��ߧ=	�L�E��u�p��-^t�Mw��f����ز�]���_G����"�E�C�Δ��7Oã��+�J��?�[�K�Y�4���xp��ٗ��[a���R#��xB�/R����I�/���L�Oa���&~ ��j Y��C_�HH��N����2b�$�oV �*3��s`�Ê�C�UW�7,�x�=��!���?���jzlx��L*ZK
�+��bv.GZ�-F��Qg�e	�oƧ+��+[b#�(�C}H���6K�)*'�gb4���CA��q�\%Pj��TE�ol�����D��(�����h������i��� �m����14QV��Ens�����à�v|ﮠ�����G1�����+�������}u5��K���ٛ��n�����&�ؓ�odu�&��2�H��%��� �!�p�.:kѰ�ܨY%�u{�3��̰e1Itl��3��k?��MTa0���. Z�n����U���p�T�=����W
Z>
�	�#�o����;-8��=��&D�(O����V�� ���ϡ��E�I$��1���CEIt�z� a�r���H�F��5br��.����Q?���
�Ec��:�<�"R�zC5Um�p�Cd-��o
��7;��k9~����6�����փ�]��r�C�`\ �'����`t%ߟXV�kUU'^-u�ΝOi�n��Yx����\DT
�dn�U�,�X��]s�FN��$��!`�;�q-➛s����_�w���mMF��տ~R�ߠ �ˊi,$��U�N����K��B�c>]  �V��E�E#�l����_��i�&�΅�8�!06��Qt������>����M��C9-�ZY2����6]��m �*������bh����,��>'�Oz���z�$�'�"��ʣͰ�:�T�r	%8�Z���ZS�W9t}��LU�k>[s��{���|Sl?7���6�xH���cS�/���6�!����<�@����©z4.�K�����"/M�.Eᵪ����L�f�V��1����$t���rr���s���1y��'�dG�Wܿ�3�ض��b�A�jn�Y
kZ�df��p�5�6���;�fɋ�>��u�x3!��d7���)uրן�kg*�����(贵�v_�p�`�s/mg�z/�WUG�[�h4�MPh�D܀�{P�7!_��O��^�?O�W'ְD�wa��u���rvy(���y���HpbV4����ן&?G߬�a�@�&e�`�W�IG�1�u)��1��,�S
�^��`+^��%i�St�<ɸ`Pe\��|Q��7p��d hj�wi?��i��@(���y�0����g�x�5�\��V12�_�Fl,svw���D�_	�s�T�"�����7%�T�VS��v�U1�e���ϝ�Z��5+�Q�01����Z�8�H��BV�I��^��M��?�K�;��Nψ� �y���6�F����p��ʜ��-�\�
R�_��b��aퟣE��d%����q0H,~�p��K,���h�ݠ�(��A�o:N\`�8��W�Z��~����՝}�yk���(a	���@�_�7�	��g;���L՜�5es����E�6?��$S��`TwIS����GW<ϗR}ő ��L&��Y�T��4���Px}�� ��,�t�����#�o!ms``����հ�Ͳ���p�u��w�2��E��I��JL�Y��g�k����K8&����H� � ok/��,X�d���M:�(|�b׏z-�WЉ�Z;��!��T��p�DqHh���Y~c��>�r�<y��r���=�}�b?�qd�YJ�n�i�x4����U�6+T�B����_�6���/����r�#�Ut#>mWOӹg7☨6�=���"���3 ĕ����s�c�}I�N�PǞ�}��Gz�� w��1�r���H+�<�,�����kP%T|��g� ��}���bfj�{�D�$}�>�7?��=V�b:�g[�h���Y*�)@�=�exr*�څx0N�7t�j:��VH�; �│���m[�_xx��sN3b�t���$�K�Y��D���p�E[�G;zJ��@��ӌ��mZF�-�/�g�X�M��Dԯ߶���z�7?;j���N��}��as��p�^>,a8�-MX�ڲQ�,��S�:�O.U�<��p���̔\!p�C���wZg����AQ�n���Ǣ��."@��o�]�t)*�p�]ғe�.-i��?%�m����5`�!��i�F2xv{��%	��M���Aū�����3q*��e�|cl1��\��]��I�x��y�w��K��H��9�m���1�r�B��:���p!b�}-�"~b3e�����C C_
�g��/�~�i���$B�1� �M<}IsP5 � cb��7V8���׸~��g?<��^A���V�/B*��V��}�q�MyIc0À�<UD56��/-ͻF�y<��n ��HI���֙��o��z4�ᵢ�y�����)��O�p��������ǜ�����9bb�7�2���׮��!��v��J���5`�$�m��L��H��������������,Hxri�u}f1��Y����0v��z������J��9����)�%t��;�J�=w�&*�G�&���9�e���I�"�)z���y�M6�I���)�+�RI��]|QF-�rjB锗W�n�TL5_1�����9mUf`P�;=��  �D��E!�w����v����W���Cf�e"�æRV> M
���8���7 �w!���O��gFw(ߠ����5f�je �O���^�u~:ףj}����ĤR�.���4�U�s8oa�̀�zѡZ(�4�i(�_*
ܳBaAl��3�3������wP&
YV	9������M�D$0w�A5N�r}�f������zj�08QWr/D�+y�/J�����>�(	=.��puMC�d��F�=�W��v�(
�������Ks�$jj�%����bt��х�/�.Xq"��AT m�,�T6'n<|n��m��$`�S���==�ᆮJؠ݄�3ѹ��ܫ P�ֳ��BSK������<��κ{.�o�����g��O�yb;!QWt/d*T~ܽ>�8{>c���WD��h
�����&������*�����'���?pd�$�:T�\�g�YD�Z;ՕO�ȹw�k>L��&�}A9��L�	 B>:CǱ��� �
��C\�v�n��t�v5�d��OKW_x�����A5������5���YR�e�ʘ�=Y��C�|��9�d���`���Nm��Z�ݎN�H�I���C���ߋ����A�F7\/E�yB�O��p�̽e�"�٭/6	�
1{��\-�1*�w�^�ۚ���k3��]�)|U���Kڐ�G���u^�2CQar�c��?:�����X�`�՗�
������8�x�]Jl���:˜3�ޯ��]��ٽ/.�/��EWD�>O�<@Ά41��5����ݹ�-+W������.��'��>&��}V�,y�'��bDO
\L�C�D���2N�CC�� �����C%���H�X��C��7/���ߌy�ZN�͈�c3�����[����d�h��Pt��jD���>&��ϢYY]^@�}��2��"�Ί��)���O7{n�d�K�����Ј�D�B�q{A7���'�� ����s�$T�;���PR[��ş/�y�Er0�x[(MY@�"�"`��YF%6�+3L(4:*����J������o�������n���?��כk-�u�_�G�@�:r��K��F��z#A
)?,�I���&��.�t̐&U?��%��3f���1fCI��^��|���C�e2o��t8��Q�s�~���d�"NrA�8�M��䷲�T��@�ϟ�١ �M�?�H} �z �g`��)���5�H��Q�o\�o4���B ��fr}���p�޹D���@�;�:Kb5�tُ/���ۯ!؀P����G������b��.)�K�u|k�U]A�+��iv�b��h0P�L�@�|�61�'���f���R�|\h���]�BޑI�0�EԷ4�'ߞ6=��zPti|��rkF�N�����W!x��00Z�KX�x�|��N �F�#7��Bt�ܔ�<�U���U�E�_/~��mvz�Uiw����µ��XnnD�+w��f��������]]��鱬����"��j�q"����Z�hd�5��\�#�#��ƿ�q�+*��D���.>�W7��Ð�,�k�JNdu�3�S�*=���U�i��ߠ�q����2e�K����^c��f��c[�I�w��ã��њ�j5+�p�@�c��'���ȱ�hӑ	W�X�\p
:4DQQ[��F�J�A(ʴ㡫`�`�;h�f�UZ�Cg6.m�m�ͧ3>�ٱL��l����/W�;Wapi"N	�l]p<e�!�堖bwa�ݓ9'AA$`i�ﺦ���o�v�L����Aet����|��+���Ԟ�4yyEӡ�l��6�Ax�OJ,&�6�z����	26�3G�Y���NRB~�iv�z��u��}+)n�CݓaDMu�Q�~%ᢣ��D��%}���ee���&V�}�?n� �*�/�N$�T���i+�\,�J�H�.2f�XO~�L�"	^�p�J���B�L�+�����w�O/����̎R]cF�N���}�2HT���8��x�g���:}�0���"�jͿ��˶���M���%�n{]�<$B��<�KK>�f)�Y�*��]Ӹ8��L�F��|,^�'��i0Y��a����ُ
z*i��-�a-���n���6�|���fa����C@f������Z�I�#���<����ebK�+�E��ؿ ��%�4e��[~����p)c��d>�s���l�mZ@ �)K�(:1 �%�%*���M0�4:����~�;b׍G�@��Q�us%��7�ಪ��y;?�8���>žk��>K4�~,��>���Y�ε��y ����"\�A�K�Y��r簾T"�D�d�+����?)
�T�����Y5�}��MY`^D&p�UW�_%�J8�ַ6��Xھ�#"� �:1�L>�#~QRs{�h��T�wXQֵ�@���ܰ��E�<�������r��Xdۦ�/��Q�o+3푆j��7�U�ZcΕ1y�@��i5��B���h�̂c�Qr������ձHE�X?�=S��F���;n�N�@2��Y ����o�\���8�qTzeׂ���uu?e�O�F;��Pz\-l�JQ��7� �O&1n��I���/~�z�bu��玛^�	B�W�(Hрa7&Z������k��?�c����؜x��C=c����|�	�l���ˬ�kCE��3�`ڼ,��/�}��iU��p�.���-�����z
���n�^������n�.��n�����.��CBi��w�����}����9s���;s߲y��X>��ȿط��ю���s�e����\�,T��P(e�T�ރ�Ŧ6��#���1H������Ħ���e���u����	�S��Qj��*�	�7��m�Ɠ�H�ե��^u\\IBhh�$(-�Aȵ�f�Q0$0Lu�J[Gb���e�(���Y�OX(wMy���C�FQ���<\j�ޫ�
������#��g9uM�2P\�7�$���l���&8��a%Ұ9G\i!���1��4=8<M��D�sG�R.$8�t�i��?O		���{�)5�A��!i!�+|cw
W(+:d~h���'̵���X����8)�]�H,��f9C�%�c�z���CF��"V���ĊەC~�E"�Q���j�Mi�B
����ZS1j
vn����&��YHL��y�H�R�#�5�������a��8�߉���l�~�+�YT�w�?�`��;�-�[ڨ�=��[H����M��	e<p�J���I\�V�T�IN��+�G�NPʏ3�_�6��ް��&�C��4����l�;�)$�@\=z�,x70�{�d�|��즨�<lyg�D�ж�����gBi%����&4t/��-�NH��i�~?���y����.�b&��Y]T W5���B{�zGL	���`T���{����F�Wخ�9{��Ӻ���t���|���{v�e��$M�4 }d$J3v#Bxn�C�i �pG�����p)���{��3a�_���.�|]T��5
*�I�{���@��!fo��p���>���l�C�_�Ptq�P�D�Y�`�a�Du��s�����8T� ��:�	h�����\> ��/P��l�xh��s�W.L��ў�j���ޕ_m��6���+Wb=�ڰ�l_,*u3��W��C��Ζ�q�:�M��W�c��\�>�	��q��H+N��7C&
�NR�Y�������()������
ҍ�� � X)����&#^����Azr_2��_M��!_�a>ሃ��k>������Q�Im	�imD�v.��:H/�Ɠ~�m�7�Ó�$�%��Y�o���(l����p�Ψ�1m1�����n�oG��$$�aK����&�ew�o3x���ʊ��FGX�:��2�(l�j���p�1C���4�&�P+�eZ6:{�vpw8�pD�
#���P�SQJx�����G���q���͓^�3��Eo,���s�Ϩ� K�&9J�04���yJ�h-�v@���P�����TCoͨr8��%�T��c�_W�Uz`���o����O6HW�+��Н/}!��7��5h���{ 7�'E?�v�F/���K���A�ra���(a�$fx`�ġӨ�C����Of~�䄧�DG�
�R��?i����p-u���G�C�"��/6�u�X�A��\�	����  ^����-��	T�v��
_p4�<yk3a�7ü2͜��:��섕�Ge�"�l���8"w2N��|�yb��e������g���2~�6αv?k1�~<�������ƀw#6�[�E� ��F��F �Eڂ=B�@���_p��\��^�ƫ�zDǺ!�fK"�\�^��/7e�vA��WzD�,:\�����C_#jk��F#	T�QX����汃H�̉�i��2�-��n�����%��<�����O�9+a�w'�߿G�Fي�%MH�_�:��*��UT�ڄn���Ʀ�e�x�LD0�?�E�����&��5����#zf1bqf�ۥC3�-v$/۷�ùW�~wbz�^��Y�~���|#���FX����oɺ��PYH��O��6��|���6�	�DnVW��!>"^��m�9/Xg��τ&d��*��FKD��G�Y�g��#E"� ����� �#Vٓ �=�{�h �����B~��GL�1�
����*& {��@ 4��B�����:%1�`���x!�	��k�~��:���,� �M��(B�������q
0�����c���]��L�ڈ�L3! � �7��׌��ЁvY��x���7G�$��dX�@����Ƙ���]	���2�C1�\ ى��i`僀|	��(`���`,����� ��kC`?���<��_�=��8 >��?rQ �HC�9�L�_3�L4���杋�� ���@�=���SDv1v2���Ձ��F��y���|��}�O���c�ՁG�z����{>LsMD8<D7�L7(ژ�<p%�,7���p�D����fi�@֩�7��\rB�;8�J���R��U6ǇX�6M��T��&����da\�PO�#A|A�A�m�Z};�$��	���Y�;�}J�O&gI�r%���yB$۷."�X�(�c]0�(v�"�3be�1��u\����P��T��$�Y����xu���(�ڍ,sM���X�b*>O�qGv 8x[PR]��f\�`)Pg��6���el�a�򠗭��Z�(*����g{*v�ct���$y�"Ui1j����H�"���zH�'���td��oHL�#䃴9��^&@9��~쿏�NC��RG=��Y8����$�@@��m�T���%0� ���$G�^0w+aC�#$������ט`�g$�L���Ag�t۱��06��^�����֩\�0�G���R��)ZfΘC�<(��}Z20���8��i	�9�ؖY �m�����7�~Z��x��ե
s42w��B&	��J�Y8�ޙ��:��F/nǬ�2~��ᩰ5�d50�Ӥ�2���S��W�d�zش_ْW�@�����9��Yz���G�T�ғuhm�a��+�6���wB��9����20
�A�� M]����Fa�X
@�~0I�{<�۴���)��|��-X��n,���߯�0	T�4i:���)Af�{��#�LZW���;�����z�;�K�Z��y�p��R��A�1O��GK���ɹ[ۨ��%eZX.�n%+D
O<�\��F ���?�'AKIɏ]Ϟ�w	�ƢN<Uj$�����F�C���������U2e�T"���5��+Čp��y@�k\<l!�mt����_[Y�c�Ld���B��RvN����Ǒ��m{��lbIJ��&�8�\j�2���	�|��R^0��B�'�JBNG���(�.���ç_��L <� ��b�R!qh_��yD��4)!�s�(����W�G������eպ��/<\
����,.$��W���
��ݍ�rI�u���c�Tn���4�����*7�]"�W�%ͳz�������gZE��� �P�&->B%��Q����Į����9�x��=�r�:��7��M��w*	�ˑ�g5R�uEy��tk��)���%�ؾ�˘�yғX�\+��Y��? ���N0
�)f~QH���.�	bs�_��Z��2�5ս7���V��výNr�Z��h}@S���ߋNe�q�6X?NmT����m��m����ѹ��_#�v�$�U� ��~��j_��H�\0��@��"<li��ț�l�n���AZ�QRJJy$�9F��Ht,�����H���o5��kfb���2W�'x��;�1=?�0�KN��+�����c��;sXWQ	G�"��4c�����
A�,۲خ߳W�9�Uq�W;s*�XA�,v�_M��i�2�_�/�[7��v�HKKW�yy�|Kx�+Ǿdm>�k�_��z�1�D�*Ll5�>C�Q=�"�D�emP.�X��]����qǥN�<��ieE��J^ş����vn��iU��}�g|�'�ڴ��	��\��KP= ���~�Hy���1om=��$V�㝟x�t��^b�a��&(Q;3�5X��6�d_���ǣ��S������a����@��գ�n���ބ�adm�#�|��PmP�n�f��T����TXu�y�u�U����_�&ݾ~r��\Y[/�~����Uj��ū<X&|k@6���3 v�ga�[O�xz���F��3����?�2���/��u�O%W�?������0ޫ�*A�u0>�H�1ޛ�%���OnS�qMfHH�(�$�k��w2��+��7��CDȤW'5�\���ޛ����ʩUg�įo`a�F1{�r���R�
���!O2���]�v�� ;�h���꣞��ХAX����5C��q�l(��8���j��6%@� �E�US5��M�R���	�]�]0���G9q�����)�=��G��C'��N��"�[�I�A?O%֭���2Н�����糍�_YPy����v|~7�Bf����,֯_�q�|��>�Lxh��l��Pm�,��Hx'}��W\|��r�=u������:*��<5}��Z=�;O���/�:��KU��g[���7\k$�o3e��X�_�(�\MS4�q����usg��M�nGG���%x7-_�]�O�U�Zĉ���v�X�Y4��-����@�Iŧ���w��o�Ec~�'�6V�E�wE+t[�P�##qJhj��^Sm��>�i�_�e���U���J�v���F;��%�����M겧�|���3��Mh��r65���v�g��4�4���vn��kIs���'噿�t�1�=�����2�xj�ٶѲ�M}@�L�+��	6�5�-c�f.m��f{��}F���'�򢜹r����z�F�~[��������g,U6'��S�H��l��Vos����%G$�6eH|�{{ζ(9qT�H�R]�i��b��YAަ����lXϤ�2I�NѶ���QӷQ�*:���n������0F2?��>�>�!��ԿY�Q����j��3I����֑����	_��댏���5�Ŧ�ٰ��f�@��j3�|͕���rX�0�3��������Z��*o�J��i������Pi��C9j�(8z��hT4-�J'%��O�,l�;��]�`�f�()�;�f��l]��������@j5�U8�w֢���}ޡ�<~H�	�T8]]�4|�1x[�ت�fp��
����m%(͌�R�vxr����_P�!+M�5k1��s���Ό�4���EcK�Ϙ����ٸ��R��>�m���6:б$�Z�� �Rz��7�v͍��8��p�]f�}wδ,F��@��T(^}�;�/q�j�O䝮�+���`�&��D�0*m՝�E�+4f=zH�\�,1e΢qG���st~^	C1�;�q���'������e#[��ơ�w�J֩�����m�p�Y�~Z�¢��O�5*�Ҷi���b�39n��\��]2!�I"��g��q�����?Ȉ Y���&�/q[1���ϣfM7��>=%�w����]����x�5d�`�3�AtC���﫷kMM�hGɑ,z�2W�辣>��!�^��*�[���&
A2�z}[HM�]�I��������h��ao��|��՛��aC�F8�����dɈ�
u=ej]&!/��I�~j~ɬ�m,�f�B�̇�8ң��Y�6<��7/�ۭZ��v`Nc�����yQ��Q`@�ڵ~G
���e,a����O���2����D�*��4���,Xw�z#_�s���ڝ��v��;=�ӶF6��-��ua+C_�� j�'6[�z���S����~�M�'���cg�Cxwoh��P���x�&S��U�\��7��Ļ�����6{��q,%�Z)���j�C1�y��&��T��&	�M��F^�r;m%��jg�O�@��D�8^7]�~�¯�������_}f]�����)XF�p�U-V+.�d�U���6�{L�WC����8��N���w;t�v�m>��s��WV�|�>�y�m�N��Hr�1��߫9`�S���U�d#��C6d25�a���`禡Jq�[��T�f�;��]WǨi���+�a��ɡ�'YY8)c����r�R�ۉyh����=���_o3bͻ�KI�#��ݿ�g����?�Y��t.n����N���0n��[\G����UC�ۄ� ���z�".&,N�"�2&%K�ޖ���G��p\O�g��흴׾�E�@�<R�վ���Iemd[�������mY1,y&<Q�{%l|�t��V����G��F����5�l7����H�7�J�GsӶC���lDkd�q��y_@���T���?b������g1D�~��6Xq�vV5�aI΃���c�������C�d��n�n➦��n�Wn�K��;���^���ܤ�9�㜏}qK.��y������x��b��j
���J�Y	����[�ͭ�2�>�BR�)��Kҋv���B$����I�k��� %����?�qЕ���^'YӘӾ�@e�KN?�#]���ڨ��R��'����ϵL��f���J�7����ܙ�Ÿ� wL�P�7� �{��C$
yLGP��1 }��

ڈF� �/
5�Y����R�j��
���EI��;��x�'̵�xO�W_5��@�K��ymn������z&ju���-�/�Y�<|TK�3.7J���Ê�Y�$���UJ������]���ى�Q�I�+�1��o�I�p�rz�Dj�n߁�����RPk��ت'x�+�\���fo�gG������[vxʴ�O�Jc��!΃��Eu����K�ndUrR�
��Y����C�h�#����樓c��ܻ�@R��%pzn/Fܶ����=�=7��� ���!�����dU��s#�=�aA�~�הå���
��_�9'�TM��vfڲH�#���\ҶŲ��gB ������
�XP�[I>����]�E~�v����;�315)�YY�R�C���x��?���a�Μ�Z����go`��TЦ"E;c}k����p��A��5�1�Q!�Di�B�u�op�8}��=^����uO*�����{.���8��$+��{?[�]��s톇o%L�ޔW��P��"a�����)-�B���]l��V|Lq�{⟤�g��V~+>=���o6:4��t
��T(������[��R{R�8��ɻ�5OZ�8f�r��7��d�W��xb�H,4���84]��ܷ�䐃!�=;�����	^o�FL�#�5xE��x!����m������]�����IGo���s���%���n�*z�F������qo��NDG� 1BG<z�skA)N���i/%�oy����:ُf�Q�׿���2Jw��m[���J>��uD9l�F��X�ٸD���I�)j�D����C��#!�_������zؖ��HB�*Z>{��9È=��A��8/j�jc�؝���H����c��,��P���A��g��j�v��
)�l,�����+&(h~��~w�����:X\�J|�$���N�l���d*�����9iV�$q�i�⓪9)�&ڵ��9�	�ߖ+�,�4�J�4,�^��u��sf~!��o{54�ƣ�dMv>�R�$�����a�@~3�A#g�Ol-�l�~�R�Xe�3I�x���s����@�M�\8�(�:���&hH������X��<��PR*`���ӧ({ *|;S�H�H#�X�7�	_ ���mS)�-�m��āg���b�"k���g��3㧣S0�m��j8���F��~Z�h�Ż���fC��3�ë�E�$���������fo.+�'s#�ȉΥ�Ѳ#�%n9���X����2#�S�O����s=�|�j���7q&$�F��6�����w�8(�;�e���e�Z���@�r)�oo�Mrko7�g�Na����_��!�G~7��{��F(�\��or�|��z�p�Ug�T��Pdq�ט˲��e�����u~��Q��ޫ{w�G|��@w�
8L��x�����B���Ƿ�͹Zt��mu�+�_6����eĄT�4��Y(�YNpHX0�\��d��N��\��"��qk�b�n������ڈ�x����/Ls�z4"x��_�Y��D�n����aj��.����Gb��(����L�["�v��c���G��K6��!H�*FIs�������������W��Dl��1 DT�����L��z�T��=_K<,Fg�e ��
�d�td3���y���W&��|��0����o���9�YǙ�fC�ȇ��-�Û"P��NG+�O�\�u�O-@*�r�v�"�⃃;de>r�k��q�i1��jI[W���(b��xE�Zf��l�g�??;zFR��'n��pt�y�z�O��=k�AGl�U)���]'X���8Q_0}g��%����n?��:c��$Fw{X���{��یVDn���)fw�>�]��;��3��Z؝W�.��I�OɋB��M	�u��:ݖ����:.��!�MBP�]P;DI��y�ʫA؛�!I�G(*��4�ȷ�2nn6�P��P����堁Gp"&f�E� �������oE��g��9U����0�����������%� �i�ȕ� dR�p0<U�/Oi���P41�����5�7[���SL©7k؀ur��Vq��h�����e���,'C$�
�qC�?>m�T�)�`
��P���fٽMsa�Y��Fq/p��Q�չ�\P�I7�@�!�#�,�Z������|�BZ�r�M}�FΞ��{Td'��!�ԙҝk!�j3��>8Q�	Bw�nq����#��v��yjpؑq �h$]/ �L	�RЛ�M���]a�c�766��-Q��#$�]Ӳ�כ���:��O�D�*=���(lU-Z��f��P�:#����6���
����w�Y�W�f������Ê��8 ��5�ݜ[���~y�&q��  ��m�P��q�R~&��/�p ��/Z�����]�4�Q�TD. ?��~jU_ۚe�gi��ݮ�Z$j�hh`~��rkG�4d�	�)n
���-��모 �w�t�r&�gqo��<�p0d��q�S��i!��g@��	/~ՓRٺ�����f���fz��$л�m�
���|�9Aշ���OO�7�O;/&�NO'��[�c��j�����ȧJ͆�Y݌iU���:WR%^����`t?����vW���@�9{׀ϥ7����~�r؛w9L$h�C���.G�Զ��翃8�t��WT��;���ά昖�Q�a�4Й?K��lji���&�vS8`��$]�^�������/�k��}Mޯ�+�}}x`6�y��]��śY�L���
y�b�4H"=wL#yq��-�����zI�����w��)j(`^%^YM�;��k?H�#`�h^ȴ��z�Q�mL6�!�ޮ�x�6���~5���n�o�>���d-WQ��@?��[��2ş�o.��c�vB�J�k���Q����g�����3Y ��&��!���+�¦⽑1!C�2�؈ٿH!�ԄQ�Q�)���&t$�q;\�Hrl�B��\��J}X�B%2�>�H.^�������M�ڃ��Pb�2��V�ـ��fYԆ�u�]�냮C"B���N�8Q�!iTu)
r�1�Ȃ���%���`�"��V��}YP�H.�ʗ��7R?�=Φ�����^~)@���)�i��	H��moy�;aW�Ν�l@�t��`H�����5�����"2$�']JE�!�c]�.���zs,ܷ-��(X�nr��+ Y��A�M MQ0�6xYM���r�5���7�3�Pfn�=��T��y1��.�7��d�:@�{h|������8O���g#ٟ]�╡&;�x�v�-���[��)��B��gRj_ޜ�i�^!/-`	���h�вe�j��J&A���3XE��%Ƈal@��H8�6��t�YJ����Y��b�f(���,{�ό�t�)���x���:�����y-�%cz��n/2J
��2���l���4�g���$�,���a�J�G���Mޔui\f�����������?�a�����97&gi:Z=՜#��
_��]�;m��ځ�[����_�V�$.k� r?����srw8���ڲb^㊚tɋ�� ��qj�^l�yڒ���>��P:J���Yo�l�?��}1^�f�s�����;��w�� �W��*��W����ï`���m�C�����j�-_�?԰a9��@������N��i#ˁӄ�.��l[�g�^��:�n/���$έ�(hJ6n��؈��v�5a}��&"�g��9Q������)N��y#��:�y���Ȫ�����z��{����fUT���l�����:���獉x�{L�ʴ�d̔��On�c���Z7���s��N��r�	��Yǆ7�pȟP�o��-S�Y��>
���Y����& w�5�Z�~qI6|�6ے��ъR'f�1�ϊB�~R}�v!3�����N�?_o|xIm
p�0!��$���	�g�\0@S(L���1	�s�{�`B��-��^�s5��GK��f�Am���+>�?{\�d:����ل}�78�E�X<B�H�U����0yE@JJZ�٬�#�̌�M���(����P������yO��y��oK�l��2�˦5�"��b�L� ���ojh�uk߭fu�Ƣ�4������J�U�k�珙�Z��M�\Q�z-6D���za�:��W�>���N�8�_a�[�����uhE�d����m �q6-��P����'�F>1m/���?���;�b�i�fy�ۀ������^�(f�� ��{��n2������0%ox]�̙�]�ޏg��`�yv�O��~�̟k��@�|�z�.9����2���U�w버�vۚF����q������+j7+Q�-`=<�:q����7�SXpd>>�H>n�Ds�
��*�}inv=�GVB~x�I�K5L��,(e�%Ԓ`X7W�*�x���ԗ�`G^���u�J�Ro�Y�H*�.�")��k�۽Wm��Z���/�vI���-o��4���ޛ��_W2Rn�E��� ��sv�����/^E-��rȅ\��4V�s���u$�q���>~���8z�[hr2V�E�]�U��N�l��癭$��c-v�R�/���Uhl��y)bxnW�n��e.���`��L@���{'���+�T��zye���:�LT�J\��]^6�&D5��
q��?*�w�R4�WmY�o��oߟ���A� �n����M^�-���7nhw!u��
�4��7"���V{x�u�����#B����1c��G�e���+�\���!�8�.�˨�����d��֦,�j��j��>d|��1�$�T������b6����k�(u0,(�/	�MB��N����T3���h�u�CB�g�˞9�B�'K��l9N�$�M����b������Z�ga���*��b�HH��4��@gͧ�ݏ��n^Ϋ$�%~��U�Ȁ�����X�4�i6?B(��Zu�8��Rw��'#��߆�L��Y�i�閍;QR�6s|�)́9$� ��B��q<_��#��|a\�#����Q	\$N��=j^����H��z�Mrˀ�y�Z�V�C��QeU�2�Sz���#"���s��i�2;�e�w��e�^��">�8h�62�̅�%X�?޼�V��Q�=]i��]o�=�S�gI�/c�oX�q"Ǻ�mr.�/�rq���>�s�ػ[9�_���)[m�rg^bURiE�Km)r�S�Jn�9f:*!2HÆyf�N�S8�X;��j�)]e�S��Hz���g�[^t�#X�tq�9�Y�q�p�s�����U��y��J2�n`j����c5e"�"�n`����>�R�����\��tg-&QՋ�6��V|����������t�b4Z�f���$�����"<8���8E�$���0�l�mڧ�#|b�*>qV/�����f����J�u���.�����D�<�7$�D��<��t6�+���T�9�8�6�'�������"�f�ń|ؿ�,ȷz'�Ũ��3#�����k"��b�%���xN����n��-�lL��&�[fg)Q��K�4tBc�ִ���{B,��5O���͟��X�6��U�-�����<������ރ,m��I4(�GX����󡤊d�-t�8&
W�o�M�y΂B_Ү��.dYZSd���d�׵����rF(3o7�����WS��x���O/˚X��ұ3�����TA��B�u�?��>�]��(0$�y:l>�	*(���v�a�t$�v}B� ��x�!�v�΀��Nm�w�7�={�}���v�n�m�	�#r#�y��`P���}&���Ԭ/����u!,HRlX?�y�h|��\�h�1�w�֍!EAN"uv���]��C�y��$r�~0z:G���<nD���|n$�CՋ�&�r�Nԝ���8��yP4��<A�❎_W苾��7��Ⱦ�����?c���gz|j���ɲ����!D�d-���.�hF��x7�󡯹GJ84uF�ɥM)Lbj�-!�B�ǈ��8V�ܿ��%3���=6�O��x3�⵿D��ў/�1�Agd�EDm�8�f�/�޾����OE5��o�}�adv�ԗ�斾��'�D�v�VɴH�"��"-��s�kܘ~x����X�#�"}d.Y�;Dx󼤕m�-�_�n�GK��x��������߶��&H�{{�4�k�j4�pr�Է�-A��>����{������oÜ���x�G��2c1����p��4�]Ь����`��]T���z��~�fQg�(e�x6�M��I�=hgH(�]�'�?f���=.�[�H�g��/�h�)�,�|1I�6�d	L��!�zt�������@��Mh��ʟc��ҵ�m[�s�SH����|��f� q�d�pU�~�w�r����w3�e��YI��R�r�=ٱDH���kC��Fl��y�w���3]���B`M�����h���#�E��H������n8��`퐲
�K�n�EU��5ii\0�$��%�Md��Ekl���!<�E��1��[޻�iB�)�e�t�}�������{S�@��0��0�d�yQj�S���䟃01��m�K��U)\sB��ŦMxBG0�1
H���&J	>�q�f[P�f1���@1QrX��2����գ��Q��O�D���s\���L!j5'�Y�D`����g� �0�8l;��
"��96�)�A�x2d:)Da��R�,c�{Q���JJJ�@�',E�$��̚$P�c��t�^��T�2�%%���c �B�sCxE7�?1������YD#PL���|���>���͠% ��'�GH!z$A��_�L \F��@q	�Å��B��,���i$�OC�� ��A l��DY��� ��1dL=v�)UȘ�a�7�Gm�cF�멂B�2&��y���<d��;��� hMA�cԐ��@O~@$���(�_ � # �2?��	� \ ��Lq�z�\l���	��-�ƀ���`˷@hH���ɮ�TK A����_�V����d���qBHH�����^�
Ї�	�U�7��� �4B�O|e���} nVA�G]".7B�&� n8E�`��-NY��9�"ȍR�jV�Y�X04�/
w�B0��C���� W��}k}���G.LKu������J��ݚJZ����\�Aue�\D;j���ҍ�n,}�He��
�su]P�����R�֒�y�z����K4D; f�hp2f�U���n�J(��t���!�ȡ�ЬGXE���a<��|>kŏW���%�Wt 8Z�� =J"�%�ݖe
�֢ʐ������@�]��z�p�}�9W�<�II{���eL�:p�)�Yc�z�)o8�PL+顇���>�ô���j���������3<�0�1X�#=��q� <���ML+�����a����ĢD�oH��F���u=���@�A���ւ�B%����p��С�N_��Q��ç~���MAe)z\H�T�Ѫ�|W��LA�2h�ܲAl0���;1�nO��%������z�0����RZ���C�d�Jf�O�[5�����.y� 0�̓������. u�OH���ej����#��J�<w��&%>X"њ�{��f�.�%A��H�׃5&$�2M�K���	M�
�#��Ats�Ε������=Е:�+�E�"D@�����YDm�����u�"}�~nyv�VZ1� �$�VLF&�2�R�6</�Ĺ��?�CaN'��}G�̈́����CH+�m�+�X�9����`��\I-���n�C?���B��p��s��Fɰ��'��������ԗ{��=��j�Ik��%3J�mw�]I�bO6���C�V��&B�� Z0��6{���|c$�4%l���=#�2	�9�F@]#,KQ4a��A�[�����x�;��Sk���䖂�Z�T5�u����[)"��2v��wA����[����?P`3J(㨈H%99Bz_��\����b�,�v"L?��D(L]$T��^H��0�a(�55�0����J�JN�8Jəz�!���Mͺ�Q�!۫u�4?�k�� F�%,���,	���/8})N�o2Wc�eպ��̷o�۪)�NK�wte������d����3��R@�i�:ޝ���z�TdrX��Z(�Bd��g��	���P޸=�:`�Y_0�!BOa��X��Hsr�z�)�u
,��(0/-)�v�z|�v��]d1�ߥg�i������ć�דɝ�
tb뜾�%�v���<����zT���PW}	�3�,�{hx/�=��$D�׼�<�z$"�Ӫ��.��`.����2�&���K���C���Nw�2�m�J+_n�%
dͽ��J�φ�)y1g�������:�m"�b'�L�pU҄���@���7��w8�� �0`P��(�����m,����>sl��;�ii�Hʭk�FKNr80ڜ3`�;{�E��s���i9��~^آ�GC9p�?�r7���#�
���I��K�i~[��4,�����0��`9}`���c���eE?�a9O#W�Y� =�f��с�-U������M��@��z�G������8���.F�?$ӿs�C�/��ԉ�6�j@�V[;�����	�A/(�O)/�B޻��+0'��u%8lG�`70vk}G
͂gi�%=��B^q<Yn�����'\Ee���םߴ�:�ۜ ������.C�^ڣ��k�tf�B���<s�n�W������ܻ[��n�͏c(�\푩{��]��zm�ٷ�6W��w{�y:���УPJJ. �����RV�g���У����̛�O�]CԳ"�vO��?���`�� �3=%I����@ޭ�D�uE&�����o\?W��=�ʳ���My�z��3����4K���g_ֿ=t��i��7��j��
v���������w��0����F�Ni9V�N�ibF7	��h�=[��~��M��z�tzZwv�����Q���dK�z(�l"`<p3�+�y2��_Z�����e�&j� �"�t�9W�\c�c���"��-�Xi�F��Vp_ֳ�\��rdL�r����;.��7�0S'�DO��E.
���EW���zsa\�����OnE��J�*#
�*8���B���DU�Ye�[Rum�FS�v;�Ы��
s۽�|�^��/�YIH+1]���5���Un'�+_/��U�	������|�K��rr��Vh1��VQ�f�D�Ƶo�6�x[︓�x��#"��5o����ѓ4��I�(�	lc�|&�����x���m�׹���c���S��8ΟK���{C�^iԹ��\a�����WN`��<|���&}��ix��(_}��*%}w�\ܳ��'X�J�h��R^�:�k�뼞�E����wk�ظU���x7��sy#�	]4.�V��t�G&�?0���㥿�7�;�8��R}<�(�&��;BMh(��A�K\Ҍ�x��B�:�5����d3Ld��U����w	^��H���>^v�v'i�}q"�sSl���Q�����t戻`��
+�����㺂��j��Dna�ͪ��D$Y�l�E�o(\&���a�\�?CJ���	+*��頱7�"~<|��:���o�'x�ƭ��ة���>?P�i�V��9��uP��ww5l ���6��"��1�r���Ź�����3�R��V��u}
��<&²(\@K�_L�>��2�I\wҶj�Ĺ�J
��#탡gSBjF�ƒ��
k���#���7�x�����FOQ���g
�?���:ck4��������Fz��o)�1;-;���*�[��?5 ���Mit\d���Ģ⇗�д��_<��+Q�ZQ64��Mւ��e�R��W�*���?^�^��DP�E",�̭.��u;���R�U��
?F�AVn4u?f�����^������>�P�_F���/��q�d�m�4�,��h��{qy�˾y�h�IP�?m~J|"y;p��$�R���F2�h���%��ػ�}����-EG� �E?��l�	���M�C��΄,yL��4�g���}��5�8�?C��.��p��٫4�mQW��,��
=	�һ6�e��H���x,g�:���.fs��@J�(���8\ǷĆT`h��n����t�w��f]��6��@�������$��,����}I,����j���66�P���k]{i�y�oI\��*&��Hd�O�Q�:&�D������7���YC(R���
Fwy���1=v4V�|˪����������i֋�Cpw'wנ	��N� ��[p]48�eC�8���w�9��StwuM�SO�T�HHĊ�IdE@H�Y,��[\�� ��o1�x�U�AxÜ$��i�݂V�%��SC�	"`t��e���9�D�x����!��F�d�������8smK�XWE����5Ua��i��Q��K�4���x��qS�Y�q󩡀�XP��Z�V>`]@}��Dx��D��v� ��l4P(po�o� �x�6ɁE�����{y�<jZ����mxR�-n����������*�rg��(��V�y^(<q���J��h��u[�,��V��ŗ_(=�hv�d���r����7�%0rW\�~��72jʱX�f� ����].*�m�2Э߉���s����:�����3��<W�#dsDX��⌬(Y}�[�6,xb�NM�%�̻첎���jyJ�]�2�iw��|l�hx�\�s�ò��b��45��9�*�p7ћ�yR��U衭��C��<&5_��)�	��x���rb���{s^�u��Y�ga�F�u[*Cr!�r��� h'tK��R*H��go�t��V�E�z�ѓF��=�7�w�R���o�UٌzL^�?��K��(n���;:�\i�4"t-�4x5֑_|��MX<�׿`Մ�}�G{"�r˶��������z��2q�^���?��f���|��G���Sr�s��&_����d�Z��2�_��]� &��w*Z�r%[s���a��(}�Z��gVF˦I��ܲ:���#�Z'>����dv�w�)��]��	�)tb�<+Րe�=�vվI���妎b���H�<v�7����/�z<:Q�?�q��M:]����u���ʴ�T��΅MR �<2v�/�J�@8��]D:�Q��%2gh�:}�,�i��9���o�/!�dwYV���^q�
�Ԋ-�m�&dl��r����뉤�*�U��6�b�M��]�y�1=�$�b����t�w��I��c�ȤR�C_�`_�ٖ�O�=yqa?޵��)�q��9����6X�|,ϸ�'0X2ϴ��H��2{�V���(��3$��s�*��/�q��#U?��@�ɋՃs�'C��/}�6���{��F�G�ۏ�\���i֡�Xb��{H����|���k%}�֝,7��`��-dI�-z'�8�:am���zE�Ǥ1�hڹ4'\7���+U^}�j�r��@*$����n$P�N�-�!p�ϩ®��l����r�Ѡ��r���@?�C�x�C{��v��K"��^G��N�WN݀�������51H�K��K�����e\i�NǺC o;�/�d�u����%/������(�r;��`���//���c�A1J��/n��P#."��h��~�H��"N4\veÆZl̘���!�� m�4,��K�j�G�iR!����۫=�'u�`'��&kt])mM�Fz��9��'W:�OB5?�����ƿ���ǘ��3.����������n*q|ij�fp�w#��*NC$�v��g�>�i�����_��<xT�t ��<K%�6��&�ƥ>FW�9 ѢЋ"�f�|Vwx�ơa�h��j����l`����[u5�<�R{3�-+������!�����)J/}���02.� �4���m��h��ލ���J�|Q�aw3�u�K���ɠ��\��կ� ّxPIG�PF�U�jd�,��rļ|��C?��í�צ�i��H����+p�џ̂�����#+T�
��N�z_���U/���#,��dQ��@��Kd��Ih��8�	��
��#w���2���H���x􍖟u�9BPCC4u����ۡ���B����1����n�{�Ȋ} �J ��L��eE�'RȖh"�/˙@owp�=��[��c]V����휾�V�R*���~��Y��S�]v��k;���e��*z��h�̞7�!&���X�Y^�	u��KP_�Y��0P�7@z��$�oC8���ғz&7RW=� �F|ƾ@�\>zq7q�J�b�dtՌ��](K�m/�����G!Z��U|�.�>��(}��~����
�)wp3H�2l��F����x>T�����5�<DJliYm�So�̭H�" ۦ:�j��t$�a���$V�Q'������|8���5���$����g����m���W3�XBlы;���O�庋�(C��H ���"�;�8������{ON�Y{��v�{�ͨ�
��P9)a �B"aO;%6ؾF�I���ʷ,�.s[��ǚBb2Q_�J �����[&���-�?=JP�/Z����o4��~_�(/����;b�L�U����I�ʝ"R�{"��d� �'ר��� �V���[e*W|P�eQ�ѩDve ��>=�!���m1��bd%R���a�����(�_ZI���?qб1E�d�.���Q��Z캨o�`NQ�NX���)A�l�w"H�Z���b��A�[��k���n�Z-��|4��
���,h��h3���&�j��|�������o��@Y�RqH�2葺�����}��`�c��-տ�Ge�n:�H����e��"�V�%J:J��B�=��i6�*"�7B�ą������6bg�6D��.��*rn��!��Х;bI!Գ�����B�X��jK3ʊ@���O,�)��/}(�7

��,�6�Za��Ҷ��7�E٭����k��Gm@\tZT�_���%F���┯��^%w�'��B���2�g�!�3���[Y5���a(1`��Ƕ��~`�uG�@���Q7!Ͻ���g"+z������F����I�?����T�P^B�G�A�W�����9����~��DcΩqB�O��z�w&:ss�d� ®z�t��3����Rm�ҽ��w�����nr��hy�"2B��Ӷ���ِtRR�mv�+�tY'�_=7L;�	vh��N��!��+�:X��'A���;���..�W(�j�5�Z1c��t��v�%�p�Ә�M��#��\@�|���/rW'��f�F,�[{�Ȳ�~���r����6Q�x윗�(�KPV�;TbJ�<$��jW�]X ֈ7�X��������,�R?N%C����E�`R
�܌���ju��	� �i�;Mo
V[�j�C��DS�@�+D �9�꿛�eN��n���q��_sI1�4+8����\��t
�x~��hyd���3�L�wE�l� S�1#q��"��������P�bd=���Q��;N1(�-�2_����b:
47��v[�;\��b�^��&�*;6]��{k^z�qл���]������{P��ǥ4)J�w܇�TS8&�ʴ����e*_O����4�N���΀%+�7z�)J��Y�ĨP �Q�X�����Y�7�c�\5d/�&9z_��b���	�of��p�O���O�9)�Id���1����(��{�ח#E��Of)F_.?���t�҅�c�"�t��{B�H�q�[�4+"#E��;���h�l-Ռ뚮��o�sM%ay�Q	�O_�~�oƄZ�
]!����!��[��z�*o�m�z����0��hL��V���_�yU9 D���ߧ�_�Ї׍���ޜL��Gα�[�>�˲o��HyC}�k}5��zuB!����rQ_�AR�wOY�26}�;�B�c)��������K,��0�3�̇���>�=��h��t�s�A����,	�u�<e"�l8��*����rP@�ظL*�y�X�,P}��mCF��^R�Y���x�j]��x>ˇ��wn%��l�ޛ�bq�4�[�����Z����~~*ri����{�7|�!�~�)�m~(���6��]�eHS�S� 4�-6�����V�E����.����5�+r��R~���1�9��lF�(Q�1��?��J� �IF�tJ�O�Jz�oO�ǡ�c7���r��P��B*��60�v��86��*`�J(�����T��y�S��@��y�m%As�i#��>��\�84z���:��ڷ̯�[����R����U�Uk+���ͫ��,`�g�"!/rF��.�u#���DYY^�?��ӱ�K�?k�� 4�D�=J�_���+�|Cy��{D9D�?��-���tQΗ���É�1������LQ�%z�K���OTWW_��tM�8�"��T��^{ۘ���ϥ�p�j���[D��y��@�_!HD=�B�ᯁ�)t��_C�V<��V{��dr�H�q���vλ<	~����epK�t0��INN/�Ȓ�{�7{d(b�}�]e��;��(�33��j�(�~2�����V�f�+rk�ާ7�'+2�����b�Ic��R..G��y�ngG"XKR75�p�ku�����&(��qSJW����ɚ�1M���Z�	���'X����{o��ߔm2�$��B��F������o_�A����x/���˟3�䥧Ӊ�>��r���@gBkΐ&���,�d~,&+xP<�5�ʹx�n������p�i܀�X�n���Yz�K')�(U0�����\�J����_�J=�Ʉ,їǕ�#�J"�N]j���L�����|����?Zdu�H*�U��{[8y`V�~
����a�y�Ƕ��(H;9�7�堣����YH�� .� ������S����ղi�W|O�8F���_l!���U�L ���b��i���b[_���Ͷtʻ�R������B%(�mn��I����c��ؚ�[,EZ����cf�>��SRRr�U�.�3q�'E>ί��=���U0��J}"��x�U\�?T�A�M��j׌����o7ye��q|�n�ئR�6��[[�|k�>���}��_�5�K�N�u�v���\V�'W)��5�x+�����^�L����:v~~�$�c�+����B�]�l�mN��}+u�wm"�n��b���qy�Gy!��o���Џ���Շ3p��8�@ɯ*P��q�@2,����f�-�݌u�� ���O���X�`]V��n��O�\��A��c�ҴV�1p��_�/G������xq��`҉��"'1J��r�~��D��C����B���)Uq!�


��?�X2����$z���^�o��"@���Z�/�>lhH"�Y��Y���x6"�y����v�W������'fi���g��m�<��S�8��7�̕�dv;/��c�����}�E6�'�@)�Uw=�;c�*�&��2����� 
��A;�nLʆ��`
�ϛh�������$TT�g�+'�*7�P�H�3����E�<0�#�'B"����=��sN4��fah�Og� ��/����c����:�;��綵�m(��梸wz����Mπ�Q��������������+rr"@��5����ɏ�b���e>����Nc����!	g�2m�:������"�J?�g�%�`�x!�A�÷821s-W��y���>Ƴ'��&�=]�:��f������'hb�l2x�FSs~x��$��V����&W:�֙$��~�E����#q��bv����x����Q>c��m69k�;?z�ld��,ž{~�L���C��)J/�v��a9]�Y��§*m�!u�z0TI$/����!����廁���"8�ը���;�$r�/�!�L��i�8҄�v�Z�!�XKk	�(���"y
l�4�����t��)J����X��P�"xo�iD��͸���h����djf����C9�.����3�}��c��j67�OJ �Z9�!	�H��,X��R������]0A�͙sjt}
K�b���L::\I�4$�*�ڒrwԛA�X�OX��z��Uâ���L9��Li^��Gg	��f�M������XŹ����CJ��ě	6Ĵ�	|:��;���� �c�oht1r����Gw�;��z�+�\�l��H$ܦ�ʬ$H6����<��Y�F�i�+{x������q�5��-�:��>M�J��	�'���Qw�"d�J_��&�����p*�6����u����W�{���)ծ�x9�-Q��U��m��o�k��#�\7]J2��hD�eD�����?��ֽ���C��X�������.���:�;l��}�dU2Ǉ[��oRA��;����\")��`��%4�B�;-�mΙw+Y��B��ze��\�p������H�c+�M���l�u"��Ȼ����w-���N�K��d�_�}k�Ά,!c��`�Q�V�KM�	g�]�.���~�^h��7V����n��z�馁f:�8���v���Z�Owr��{d{�J����Mƕ�G5�����6�s#�U����D�������8�k��8&�p�KWzcޔ�f/��\*[*.ʺԅF6U���ɛ�]�7���u�VD4
O��3���0v�]dh�g�|B׍D�c&�pv�M��đ�u��8@\A��Mb��S$Q��th��AJk���b�E�{�5�2�]����0DZ7�|������z���ߏ(�¶r�D�7��!0���F.���bs�8A��#ѯ��_��
�x��p&V��0�ND"QD���N#�ۏZ"�ʋL(ڷՏ9!V������$�@�q�<bһ�.�_�;R�l�$n���Է��qbuqq�`|z>��a/"��$�p{��#�1H���?��mp}��������v84 ��u5˚�OSiG]����_��eR��;��Y�X0oM��*�6>�U;�뷁��e��b��J���-�k�Zڶ Y,^y���ɫ�A��yL� ���_�߮��vbu;t��,�ݬN}Y������K���ak]�F����fj�A��Q��Nv?�ޓ���_(캗_��+��dmt��b����)>�~�$.r輫*��z]݉������)aˉ�X�)Z�ɣ�s�dc��E��5è�\��?QVģ<��-%�RsM��*^ybȸ9e��U�ü6W�c�D�w������<c���ڄ�$T��������s��C��!�� O�7�y�(m������ZX9k�>���v~�P<:�Vz�B��Z6�r�ȍ��~1". U�M�d19�l���\l7�KRn;�:�f����O'��9%:�&=�;[Y��vd��{n��~$®���x;	s���7q`��؉V��0Q�m�gu�^���?1�5h�ʢa�_��։�Ly�9;ǰ���!����i���^}h�pq2,m"�ɮ7���+������Epں�e�"܀��j{�PC���J>�oz�0X��]8������R�|J��n+r4��F��b>�qgk���k����Ã���@�|�Lx�PB
�wv�iQ�F&D�!p����L��t��U��i�U~h,'@���4��)�x�A�G��E������UV�{9җ��H�~����u�$@ko14�!jY_a�p��ZI*l!־�D��ؠ/f��� �Wg�V"���`�/��j�kz��`�a���
�G�s0p���'â�řR��o"�{��I��)�؇ u�_�Vt=c���?��2߂1��F�D�;&$C���䴻B���(�9�n&)�xs�#9�����?{Oh="_`9f��{"�=E򕇝)g	&������q�|[���{B�wo�/��2�Tžz���< �VF�$�5�.��a|�%e�q�,��Б�i�iB��Z6���5(YKV�����U�׹(À��,�xP+���Z	�q��g���d���T��T2��� �P��X�Tl�Qh�S��%l#�vZ
�u��h*�Jb��X��i~�T��)��G�����{��ϗ�Ϻ#�3�y��*V�ޮo>��T?�p�;��B�q�U�)Y*����9A�����	Ů(dL|��Sr�[���A�G�⛀��&�/���7:��	�*�34��G��*��L�d2���dɘ��p|���ld����Z��{��i�e,���C�2��@<"2T���/XA-_IB"]��k:	��,��)L�&��
�`�$FF2r60\ƄΓ��Kg�O"c_5D�� T��,�ʩu��*Б���E���h,蚜��yp�Xa
1�І�(^:l�f�J�0�L� b��"0�%L9o9 ]1��	��}�9���
tM]蚭�yBp�Ԡ���������[�	���*�Ua�:ѯ���F��D���7�-t�tm��C}`Cx�5�`��-j�E%��HǀjD�Hf�\آY�2��U�#��g�NK�CǦ�G��( f"Oؚ��#qÄv0!t���1��U
�֚*4D��/�*ĀY^U��Y�(��ǍT��b�B k5.\�'845��kvLv��W>����}���Մ�°Vl\NN���x�̆�!Z{�86�Pl,)�e9><��"�"h���p��#D�>��/���uR���Lv��?�Ċm�ɚ�,��JDφ�;���~+��=:>��_���N�*���?T*Ygr}?i��{�E��vme�:T�L��Ǝ/��a��U	��?������P��k��h�P�8T����Ăr>��b��p�T4N�"Ƥ�q~��7Xj%��Hx��%�퐙@�՚k������'vBK�R��6{\��I��q�H�lh�=xı��E4M�+䉛4�,yÝ�
n�#{��"�1��ό�9R)�\��X �j>��i�F0.��9�$J�S:�m��.��n�)�@�}�N�\�ԗV��J1��	)�N ����:K ���s�	]~��/�Jk7�t*�<�
!RBQܲ ��uvb �����;����OLF")�S�M��$��U�,=(�i�_�`�%W�+� �سy���Xٚ~{~�,�vI�<�=@�.⊆	��)���ЯLC�~qi��ǡ�C ����p�K��i���W�)��;���<��8['����C��%t��N-��zMm#��϶Q��MH��2��T<�α�И��Hs�}�	;8q9w�~����ާ<v�����QW�@(�N�w�<M�	Z@����!��l�_�@ri2x(��H�L��ڨ�$$[/��cg��	=��'| �͗����]���8�}�d���y���&>�!F�)�NN'Ԟ ��î��G�R�~�z֘"N:6���6>X�����v�:}
K��������*�D��Bʙƞ�^_��Cz�>�q~���䙄�^��>�ʵ�_Ez� ���z� �P?,2�{O�_혭������70���	7���ށͲ	ox(��;~�� �ꨥ�FQ$Ik��9�~�Җ����% ���;(�a=�Ҽ��0�ɍ�M�����u�[x��<f��])(~�rM*Ǹ�W�2M@��S�G���}P�L�o�+,w%�mu�^
�:c�4��ဏ�?tx�P�J0�v�_v�GD��;���7�x̎]�=�=�>H���[ͺJ�m��
Q��e`!�|�쌍W��H���F��B8�n�Ф�74+m�Y,�'}Z�70
$�6��O�C[�ͤ��r<���A����]�o�9��m��՘'����4�5$j�<�JE��c[J5�M9�oId~b Q���QE�֜]̈́�~-��o��\T]�6�1͕Z[q�b�$�"�=�rw�%"o��P�d]=�עr�~jv]7�i��3Ncr�ӡ&`?2��;�d����h��*W M��a�,Ǩ��om-� �m]��N�!� ;��=��£ܮP�h���� x�p��b�߁��j+��C��+�	�{nP�}(?�Wc��(�e�ɈEL��~��C����1����v��Sf��;u,x��Q?�/�]Q��r�GFPEQ��4R�	5"��	��-�?5TlP������#�G`A�|� 1��P?�w��&o�����@��4�&�5��w����d���K���7�]r��C��?n��w@y=mN'�`o�F��I2ॺv��d�ȁ�O-��\�!,`�GΆ
��v2�㈡�@KE��F���J(B[�\>cTi�R7PR�M��b�U1��bj
]..+�o���Ϸe�W�����z�?YA�Q��i۱��E.�\���1�����G5�+��f$��p�������m�b�����:'���~%%0�Gc��m'|���?W�BL��ʥ����9�v��;�l]���q޷������~�ތ?NO���V�Cى�|�{Z#�e�*{!g&`-u��SI�}M�[�����p	(��d:�wVds�C��%�s��QT;�>H�o������ �^�A���&%��{u5:�LD�)W��Q�K��i�1;���yV-w��&����|�j��J�%��fcM�A(�W/��A&!74��L���޿J�m��^�2�ͳhǢ�O~���{[�(��f�0�.k���ez������e�+�Q��
���Ϫ8���+Ø�G�MNn�Cdyo "�-o�b�ܰuI���u��"L	>s�pI��R6�6��!T-�r'��G�(��ZQ�%3	�vi�li�~|���/v����~I.�*<�r6X�+�s���,Y�v�cȘj%�7g�*"��CG�#��(����@����-�jq�X�ޛң���-���ȷ�.%6���n'P����я~�$�,yM�}�X@� z�s��k?�-C&{ �^QÚb����`wn�|�QN��o߉�u�$�T5�IY"�Q���Mc�}o�W[�`�?��ސm%����h�-�]��hdEt��~K�$��vx��+֎�w+�ް��4��tJ�+��Str���t�F�y�q���C#6rT�@�J�ş$��mΣ�6��>�L�S�D��Q@��9�U�$@�-�v�cJC,*u���fۧg3
�(��;�.Ń>��z���$�x�gW���[9Ky��1f��o�{���b~����;��%	��X=���Ka<N��D�.h��#���y�ļ����^�I���g�ׅ��*�@�_äg�I��`D��k'OZT	�@�t�rSaSX�;ė�<@���$g�"����C?~�5&��ڣ��V<%��e+��̳.��P#xY��F��(�_�˰�uBFi��j6B�?�6��'�?@
�����91���Q?(_��x^�S�I��:��b%_����;�6Xٲ_I�z�֢���~�w7�����r���~��5�K����}$*$��>�D�ǽ6z&7� ݙ���(e�~�b�M�)�����?��Xi��-��R����	�ݱ�5K5��*=�~��DdCV����1�9�a�f_�[
���4醗}΋d������h��,�Ơ5�"鍻'��X��������.�DG'R["�aҰ]���P�JF�^�Z�׆�З6��5�jrW`%�#h͒m2w6;��+0��<�	Ѵ�k��|�<9>��H#�hi�ٻ�@�{9e#���z��%T�����4K"��hn6���#���t�� ���ӓz!qPNy>z�'Ⴤ�VR�}6�!s����j,;�Xa�wZ2"eqH�R�SJ���Go�	}͉n�������))h{����k2���Ȱ��.{�'�峨��j����C�ى�r�o.G\��I�8��,�^���	I�o�?>e��ڹ_g�}3�ew�����p}=��i�w=�XJA}�iK���=!]�
��6TO����e��e���p_�yz��?���p��� l�m��N��|ο%���3��U�����Z�n3F/�Qy٫�.a��Uki=�+Ccp����	�*D���	T���R����	�I�F>[��OF�����:S� �#	IRj~��f�Hn���UAm�G�r֜�clT��Ɣ���7U$�sא�l���ܾ�r�Sk�$���� ���M;`�N����J���%�w!H��'}��(-��L �f�yG���}UTR��Y��r�h�������C]��V��)bA��
Ηy��Do��(�a5:�_牤Ə�|����L{�c�z���h B��Jv`�E��Õwv�(O8!��6��S�>���0�F��T�P%�w����>�TH���.��*_�����}�����fZ��Y몬۴i=��y�$�-����� e%%W�{/��Mw�N�������������$����6��K��"��%�U�TD[�M�~_�QIΫ�(,��m�冱����T*���ŵBq�A+�%ǑZ�g�sF�v��"������h�_�X@(���[�vj�|y���uH'}��E��{-�zv��]�q� �������_ח�4گ,�1�����@�{v��K���D ���/�Y����A������x�l�oF�����3lE1G"�t��C���%�/�k�Õ] Xכ�'p��?�忤����/|�yڃ.�8�lĨ6��).�#!�p)&-�`<�cS�&h��r�*�3m�ʵ������D��WD�1:��`����[[�̟=��-��Q�)�p�����Kbrq�!F��>�m��(>|?!%'��B��(��b����>7v$�B�3Yu�����Ž�ǘ��F�n�U�Q:Z�{��fM���6���W�y�0���u���{���ұ#�������{��w��B�Irj���Ht�Q,]�x��AE��9����?d̈́�h��s�@S$\i���P����C�g�Y���K��~�=;-y��u1��^�~{
�2D@���4{\�|��x��Nl���3�u�:Z������"M�h������̷Qև8V���C�ҥ�3�����N8�{�L��2�G���*p}#��S��|cmٕ�oS`O�1��Q��l�6�R��A,-�
�:��{����+'�!��~�3�4�W��/bf�*( ��Ջ���$��V��[O�i��Z<b�*B���r��6�᥆�+��7Û,I�cbb�oI��߈l� ����g��m'^FO���oty����ˍ5i�s��$7�3��JFX�l!�쪹&�A-��-�p_��:�y�d��hE/�V�f��VCx�����2����4	ȫKƸ�9aUD�U�mRi;|��Iji��}���o�XaoINq����'t�*�	!��I���	2��Y(��U�w�3^��=n��y���;�X�GW��i�?��֦�B��z�J�>��9@z�~�y�����׿���s��N%8TZpLhrS�n�7ם~��7w^�Jbnf+��f��f��˥5���"�qk���"md�(�VKeнф5/ԗ:?���G��M H�\׷�O{�B��o'6v�ǢCVZō1�#�.�O<l�8�9������
�'���wD�O�T����m�G������#�XD��m/���垆�Ӎ�����Ƞ�~d�	!�^��}>D��K����m�Qq�1�Į��K�6���AD�Y��}��'v�m�'˝�/SE��M�Hi��S���!���{'{�L��7��r/����r��7���׫����#�	��0s%jD�O'��1\)�Vfj��&��9� ?�o�/�wS�c����g&B_����&�;J�^������|
���G����ή�>XS����g.��2���|�GJH/�e��CJY#ğ3&y���Y�IzR�������1�ػ#���E-���a6#�,�拾�0zU�0�� 3���X~��s��O�2�I�� �!�O�|n@̢�����Ɂ��?�=�����r�p���+��H�U؂�-&��!l�.�j	�o��H��~cƟ1�'�i2�-T&d4�4ӷ�Ѥ�R���ƭ=��������]��E@X��2Fn�V���VІ������i�Vv\�x)n�ζ���g}`���p��{�bחʶ������HA�35~�E���dD�]��R�#� .��aa&���Ɠ$��!�c�h]*"��EJ�[Z���ׄ�lK�57�݊3�Ņ_�hDXPII���{U7>=�ou��/�+�LLVjӉhԬE>�����R��x��\>,Ҭݨ���A7�����E����8̛�Re��1��\~�W�U�\�a�
��^o�ri(p�_ř(jݜ��/~]4>��;�BS�z���(�I���W��S=Z'�r�kQd�uhE�l�M��j��>�Q�&|�_����l��,�s����"��v/8�no��I�E�W[�]�Mq�˄*0���v��v���eһ�}K!�we��Q�I3�E�1�W��%D���/5S<���k�o�H��#zi�(�Jʎ.��u�'�W�/@�6�jq!-93����������G��Gn��D̘�6rE*Wtj#5�`d�OE���P�/�� �����	U(��BRv���Ф<�+�e$	w}϶�IUGHSO�K �ʐo &�Fal�0��{��d1n���/}����C�#3j�3B�q�Y�"�YhP���4p��ګ5���D�c`�훏T��eچ&k�]礜��wa!���^���4�+E]kj_�M�.$�8�☊j��ybm��4e�e��o�����c_v/|5�)��M5����~�]A�����M��r���}�M�ܹ�eA�>���Y�MB�{��!�8����sh�˕u��2�<I�/%W��P�^�:d�#� s�H�,8����)@��g���r�q����c��
-�A8?�#��5(�O�U~4B��p�i/�-�C��焤;�5o7Y(.��eXc�1vޟ��x��Pa��'��4��%�y�0��Q�����bFkS{����i�2Ϫ+˦��Ĩp�g ��])�t[���!������H�)��� Ԁ�yI��N���ǒ�Ui���u8R�X�����n}���S�DŤ�L3�f5��wX8��_{~�G'�0�s)��|�% b(PoJW1Fj�_8��=�d���0�Iu���ݚ�H��)��Ϝ��wP,76�]�?n��N^,<"#Q�7�4����+�岅J,j��nl����U&����$�=a��\%%)>�'�d�KG�{S��$���ʌ*�$[M_W��[0f�T��WC�P'�!]g��mi"����[H�~7b�0�����5q���}C�7s=�Ֆ�ڟy�Dն��]#�"3�""��p�7��b%
G�l���RM�6���{���Y�O�=>��u�9�+�1�����aAQfJ��aJ�����_ ZEF�ד��.!��K���/��r��O����U.�NqI��6�;�t;�땻��%c�0��>̝�2�2<Cݨ�G1���јS��C�<5�E�(Ig���;f�JLW��[4�+����#=�p�j^tۊ3�� ��D����/��`	v�W����;�Ş��x0)��4/��B�\�.�4��_�&@�-�p	�ػd4���m��u�C���5Dz��tŔ?T��g�[J���Z����[*��ؾkM+.}���_���$��[̆m�|~�H�(�B��{Thvx/��IQ�r�~��[[��-q��n:�$�N�Q7���6�� i�3�#��fȜD�S<��Νy)�:�<&��M���s���zgtV�V�2������U3G��cJ}�������b�fiB.�w�����_5��O�`* �!D��j%�4��1$�3��0#ѝ������*os���e�;��a$��6AԊ�:��w�bB�W��zlj����0tF�4�J��(V~k��-��T�_�]�'�ͦ��G�-OfIeDT���\L��k[)�����^~��.g>L��Q�ةaˌ�g)M6����\%dnH�9В��e�I���G!��	��(� ���Ou�{���l_��Z�_�S!C@��u����:�Ϲ>�r�
��-���O*)��.�ֽIO�i�p�q�$��˾���,�XsZx�Г"L|E�������à��y7��'o*�5s�Sf�V/�Fy�9q�t3��?��	�%�?}	�=�����z �����������gR᫅��eq���͍|/VĠy�:�3/ �cz>P��_�p_v-�L����|��o����Y6,-��&j�8+ve��B�i��#q�@�i��]?{ �a�[���e~E �u�(RW9I�Wʤa.�Ĉ�:O1�li$��&��(a���J�����ٖ�	m\�$��<$@f	Οm[&�;b�换j����B�/���ET����z��pB�|Y��� ���X�l��k����'��[�H�ou�>�,�ON���'�8,[֐��Dg�V6D4h����V�1�\K��q��g'坮����W��'�|\����|X�	o���j6V0ii��Bk�������Mc:�z�%jKm���2U�tt�%����3��[up7~����(�Т!�QY3Z@�S<C���;��.�\�s+ծ"��[�)m�:V͛#|˕Z�ˈ�D�@>a���n<���੧jv���-���O6nS+�#ф�׽ ���?���g�0��,|�.nc0V�)�~(��t�P����vpk:)��tIԞ;��C���yK��$�bI�%�������)����5���-"���g����9�`���v1}��'Sڅ�`�ؽAW���� �z?�.����o�� Q2<y��
���$��'QI�ŒL��w/�7�^���GsD=
-��p��o�3��>W��J�#�^5�s��A(��@PȆ�P���F}�ˏ��l%��v#����a� ��R �$����}�2��ccn�=��82����^mu��p(�w)Z\�;��ww+���Nq����;��������Z7Y'�I�ܙ={�3�K)A}N���?1��h)D���x��Ev��a�0��X3lΟ=߀�[�����Â6Zr%Ybv|�=v."os;6ːs��8.B�3~b،cT��n�τL6�H#�e�[���'«q#�|�NkSA�XE6��zl%=���b!3h"\C��{6�'�z�In$Z�%����zt�;��t��o߽8��y��*��䞷*!�X�ٱ�*�Koż'�����b���)�P�
ee!=[�1�8��-����z{{C(�^����M����ި�~��\�br�j�t�sN�-I��`�����e��x��ȓ/����OT9�z@D?w��|9f�}���km��p���L�,-����	��Q���]�N({�*^�����Ći��9l���v�P���6�n��m��Mz	�N���H�镅���#�-GV����
ѻ��1	����[�0V�� ͷ�]<�y�0S5���ɂ���?��0Lo�ݿ���,'�#��v�Z�������[��Yb���<�%gZ:��H9�bl0{k���K����j�iS�+��E1v�����]�q����L/Z9����4(�}���!O]�|��o�}�'�� jgԆO7�)Xک�l��i�?*{��9�6x���
��E�Ĺi!�r�-��??�nsB�.7�&�M�D�Fl2P>�p8��j;�V�Y�.YBkJp��.E�]���	ҏ�Ԡ�G�hUqGk�\yt�s�-�>v0f	�B��֖��ꆸy�u�.�r�,
;��:�$�}>F.��@� �c2Tc��S��Ni)9A���H��z_o(�:= r�|P؛?λ�jLpi�t�y�^NT���n7�T���M�K�e���M-�>P��9+6�P�?g���K��g'C��ٺ�F���o�$>2;r"W��W�k��	��݈`���`�L�y	�P�j?��T�9v�k�֏-\<�"��ڨ=L3_���y���[�!��SG${�"�ɯJ����v�#^5]��5���&D�U<����i�r;V`�s�
��{G���
����0����ބ��L�g����|�2Q�v�����}��_�炃=l��>Gw@��X᏶�C�{�݋p#��m��;fy0�>יw�&O\Rj:=�0ȷ�u�~ϱ��3�4�̕+{�t9�i'��)d�v�P���V���*��ظ�̔T������D�eP��F#7�]�>���Ǎ�Dԡ�ғӁ͘�����'}��2�r�2LG����j����1i�V�?"ѫ ���g^+��{3S�x�M:�S�ܡ�c���n�Nݖuۏ�(*cy�+:9h��{�d:��Yh�@�Z�f�Ew�$�^L�tԜ]�XX0h]���SL`mOB��Cr*#�hbӏ�-�w۾���nQ^�f���J�{1>+8��T��ZZ� ��Xs��c�{f����X��7�9U�cC����Z��Z��4�URq��eS!]4Z�y�eC|��R��� `�%�Ƹl��^Qg�m9����T��	&<�&��[�o��`���DfL�;MK>��n���g������V�bv�y������P;S�]�jED�p�z�&7�_X�6P�1�;U"4�[&-G���Ӯ㺰scN��{�YV�Hj�FP�;�+76��kw~C�^�ɍ�V3��p^� ͕3�?����i�O-���Wh]F~��[�@�<��^�zG3?����Z0#Fn�ܮE��<EJ�V2�bs<Q.���rV��f3�"�L���h��1C��)�oo�{�3:A-��z|��JutR�cpd9��7T������]�ϫČp[�`�Z�_޴�;��x�wϯ�=�WV��r��L�1t�Rg��3��	xd����^�\�E�CH"K�z��=Ҋ�DHI�����d3>Xә�PѨμ�yf�_�16~#F=V��/P��0�Y��Rjؑ��d�ӳm���y��ˤ����O��C��O�O�c%�3�o��iz�k/r؈x��%���SY��v��̔=��K���o���O8j�FN���fi�Rᩂ!6x�R�us��\��l����w�\d�4����UT[׭3s~҇n�ŗ\|�?�E�,9w��/�C��h.�����A����e�fb���$F��֌_�Ɋ�|41�+%�����::o	�K�����jB��_&)j@m�e�v\���x��_�@������0�y���g �J�b�lٙ�Qb��e|�bTО5���J�H�g������0�x�w�D��<?m�N�yЉ��ӄ0l����F�����1��5���=�@u'a��(.�*�x�6���_)q��͛�J��j���[���4pbBZ�����G� ���d���f�v���dN��\}�("b����Dq�4�`��7C)2H��Pغ�����'ע�ƕm�\�c�;p�%*S���?�:އ���ο�ij�㘈�������Dӻ�����`�Av^U�����y�Q�3���"P�k9�^vG��@37���E � |ئ��v<J�e!�F\�W�2  ���	P���h�U�u\]�v,d� 9����j�3�|����6��/w݆GK�������R���3�#(|W�6l�]�#Dm�C����L.&��>�q*�?� 't�}VRB1v�oɓQrѻ��>cyz�.�v�^Ptu2�F����~�����h�G����~�����L�^M��F���F)��8�? ����ظ�災#,��A|<П(���PV1@Jf����? ��@���ʘ�?���%6��]��48�������0���$�I9��)����vﲇ<Nd�C@�0`6��$&��y�[FQ�f�����c%;���ֈ���@�Q��a�=2O�k����%��N��OҠ�~f��%`U����w�i�_����{+�j嬎������܊CC"��'62�\Lv
�iSF�U<4q,}�?��'��B�`�Զ�ZO�/'?�@���j����hh�v��rh2<���N�e�z0ꓒ�nTn��s��~��G�t(k4��)S�R]����t?q<���o#U�b1I}u���u2��87��8`��1���S����+�,zv��`SZ�5����2��c	��B/d`4
��퐷�/^�H�0
�7��[�k��,Ab�`&��C�с�i	�=}$��n^���d�~��B��������*�����^���	4P�fI�D��}B����"j�Q�,�1�5�"b3�,���Ql��/P\4D"7ȼ��OT�������uǄ���I:�-���X.4t��L�7�*�g�j�Cq��f`A���(���@����*]+�����D2�O� ��$�a�ָ�R��@�"��#P���b�d� ��I�:�ݮG��ɱ��\;�ܹ�\_/��V��x�6ٕ��1Y�x�?��g�֜%BtF,�g"u��_�8g��q�(j��u��Qjd��-u���6��Z�R�#Ip!��(jE�ǃE
S��p�E�m�vb�\E�!� E6L.�����`��_�4���d��E/�Q��.�,�H�4�n��!&�|Swsc�yV����֎��k�&t��hi1dT(<;$zL���j�ͧoa���]��Mg==�����~V�M�W��"/�m��
V9��1�	w���4��9EP��C���ÑaC������k���a���%b���Z�
����������,�!��EaJ�_+���7?Z�{�S,>�}�^a�k�80��ml����O#�b�⿏��p���JI���o�@H�YHrr�_[��J�	#�����$�=�޿�)���>���gP�tЂ)N�����͟����l�������Et���� bӵ�mp$T9��{��)U�X�ʮ�`��g;�L�VA�Ҫ�Z�!	�Ղr���V����`1:�p"!n�
O1�aYmu&��f|HW)	2�d67��V�]`�U�Q�A��ڊG3!! ,Z���V���G��Ǯ�'j�����m�ڑ/=9;/���V���R�瞯8\Wk�P���>\.1k��Ng��f��a_W�J𳮢�p��Б�	���`��/Ɍ�\�&X�L(fA���%�����WNc&H�tC���i��!2���Z��r�Z��Y��=�l��.�\�+��-��$ґ��6�_��������b�R�;ʾ�^'������*b�#~��9��`����g}���V���HF9.d�����4}��[mgqtt�Q��?�9��ɼ/(赵����j���.��ʌ_�mİrZI�4�>��;����<_���@E[n�ڶc�m�
ϳ�f`��p�F��~�3[]�=m��[�d�"1c�;�t��l�����c0���������^����/Om;%]LC�j,�)O�����z����Ԣ�#m+�<}n�]e�ބLr@��Pf?��l�U|�<��1����P7�}c)��O���C�5ttI�na	�.����Yr3et5i9�o����'=:Nb�����s�3���'0��^F�^D�J&�E�{��K�6���[�OV�\�������P�Hez!��*Q��'�\���P_k����ls�o/Pb��͎j9�E�S��w�Ck���=����٣�C �iy��f	`�pP�p4FJ����lU�������7�g�r��L?��2g���������p��*)��R�)fAV��8��Fm���ݍę�t�ޚ���!�'rc��8�y�k��Yw`o�[8LC�)N�[���� �.j�]h��)�\���'p?�`��A����B�%y$�����g�����cT3ɒ��*��d�Òk�ˍ�1U��xl^�b��"M�r�Z���z)S];�$���}|��1�%��GY�XE*TH�I�I�z��N�w��I,y<�6�c�j��W�b� �*�x!�C0ʦ<��$�f�3�������z�xVC!��rЈ��0����$�;��͛$�50�ǋ6u	6��"K�l�梍 Z��f�^hF���\�{�݇���J�
W$�p�Fܿ�j�3�9�O�v
<h��5;�^l6�jG=�#�đ����~F�R�]�
���?�͓�(��w�yL(NY��{H�b0l�2�!�!��
Ж�]YAr�ǒ��(vG�s����}'���/Ex}�r�HTU���q^�{��[�"c���'�?P��;f�/�SY�_�����лv�t`�j�4ج9����+U%�,vȀwrd��Z
�~���h�H�>e+�� 7�t�h$�.!73�}����ľ�"��q�xí#1]�������Y���u�������۴j�C�!�~�������屇���r!�9�7YV2��p�M�T��/�"��yն��8�Efn�>E���2�1n��� �9Z��?��v��U������?�Yv����Ax��G�x?��.�6g�21,�bi�e�N��B��T��:٬���R%F*���9˝՘�G�d'A��dH,���dS�c�)�N��N�Jݮ�����B��?���6S�6R1�"t#I*u�<�a;5�,=�h��Ѝ���
>!u�z�Hȣ�2T��ڊ�p����]�\�}��\*���jSܴ��� բ��Jv�54�(��ڔ3�Z{03���8��	�~���#���N��V_��r�ӂv�� (@=�������n�{�a�|�$��t"8c��3"Dָ�-{8*��u�<�/2�(B0d	z+�y��Cn11��9�G���uؤ�f�Mˊq󐺀���о��L>�#u~g�5��'����m���:4��G��m0Y��k�_�_���<O���j��ck:� �9�fΝ ����]�!���0�~�l��u��m�&�
'F		hT���?=l�J�O	4p1D5�g�^�M,��m����łK9(����G�*X�!r���Z�zަ�c3X� px�� M���������G6���t�~/�Ux�빗�D�õ_<��c���}��*�f���o�����V�!d�:k���#=��b���⬽d��}qwG�?��q���z�=7�\s���pa>���yic��2���}o��k]����<M���E^G�$���l$_hp�?�äa!�x������`�M�,hm�=�G?\�	���|3{��A���i�#�0î�����q��Q)R1��HG�	F�g�k�]�oÚkٳ!J�F|LF2��l�Y����f���K�)?��v��	M�1V�;��7��XhYo�mP=�i�۬=hXC���$`
�(���	��~.0e�2S1h������";�Q_-�	�4T��}��b�\[$R0��H)�.kB��V�j�3�jeU�b��T�ɍ;��Pg�4mC�"�_��x=o��:k�"D(ɶ,/���Zѕ8JY�4W��\���� �6�����y��v*�����L�
 �r�k�������?�:Q�mL��w�R���HH�\��K�]��1o5&%[����D���~&V�������h�f��΃�i�йSn˄��g����}�e6�Y���ˁ����l���k��0�q�d�ď�:ÿ�t<Xz`螏�i���U'K�~�����ss���R�Q0�,�8�d�FҦ�����gw�Z}��Ai�٢SkQy6`��̻�8�ٻ&E$ɱ�[�q�V�!��q�� 4\�f�v+�@]���_�*�;��b��&�3I�rw�^8%��r*{��it9�o��0�����-m[M���w;�?g�Kψ���6B��BUZ��bd�	H��yc�s��*�?�.�}.�_^bT!��
�2���:^��s�Bl�r�� ¢>�\f�]�k���,���Y�&E5r�"������1��b��b��P���z\=�ծ>鳸�X���Uh]��f� ��qxx�b D�i�%�elDA�[��!�����!��i�|¤e�s�4f��XD\<^:	چL�B7�bd��֦m(H��ܙ���n�v����������vi��o��Pa/b�'�zI�s�B'w~.���t�o�,)/M!>���pIUS�יnv/3O�S4x��$����	I�ts��g�;o99]�*����۩��uIOCH��m�o�8rW3��-/N��D�L�~7��������l|S�ũ
s��]�7L���! � k���� ֵ����ID I���g�Q9�P��˿7X�;`�;G�{���O3�L�_��џ5��%���P=�[�rq�;��l�<OĜ�t!�Ћf��ٲ�S=�|5��qcA�Z`�KXD:í�1F0>T%���4똯�6�8�7��P�2M�����.FT�y|�����`3A�]M��KpX6b�6tC���u�dH���;K��9��������(x���M�����B"x=��I�Pl�;p��\ �L~�X���^�KΘŭ�%]��1g=�緍4r��rjѝ���g��9����E�GZ햁���L�� Ka!��Z��p:��ߍb)��������DG8���fg:˦"�>7��k���r�P���K	8f��{8\�^S���f�W�,�x�K˭P���H	�@5��9[q�]��%"��E�'w�V�X�o��D[w�nҨ��h�ݹ�LdzC�����Oj��|;�X���A�c��Dm�e�[�|�j�$�TCE�4�� �c�&�f�L�@��i]^G�{�C
�뿸�W<_J�#�dK�g�5/g��/b�&���VP* yC��;�l�HA`��S@1=�ՆL�e�gc7��v>��`{N[�a����jX��M�{�+�2�8�dg���-Q���)_�����W�zb�e��,�����:�r^�5���;�
C�?��ϰ$���4eQ'K���c�_�*��K�	�G!
�����ô��P	g�S�j������
�A���5E��B��;�L�7fH>1��؍�%O����˰���zSPg���&���ET/���p��E#�u�N����Q�&&P�I��)�O1^����V|䳡�e��muq�Уq��R�0��ʰ��+��ҥ�)`�]Ğj�bO���f�6�N~�f�u�`��ui�w�A�����A��m�6�CH@R:O|��_�Kk(M�k�ά�zRv!��pd��~`�~Sj�'C���Mq��Yj|�<��	��5��9 �m^Q\�LbwvGm�}m"�,_V�`��~�9�����rA���P���Y!HqM�L�.��b�g�j�P�:��L���NsV���:�R�}�Ψ�fe~n_����X��̣�z2����@s���	��k�N+��y�����M*(Z���tN��m�?��y�~1fd0H�^���^�Ikm9��1�=���1��g]��%��j�-�SY���ę0��,{��1W�3�C��
|E��s`����9=��~5��&����T��)�����v�L�r8�MB
�U��#�~���."�.��2��4����G�><�A'��p�����DC+R6�$p� i�~).���Y�'K��H�'V��v: �>�����u��@pr�.�T����&�Ўg�nA�qs}���u�,2��q�1it
Պ�ȥ�2�/jcq��hy�$~��9���@�G�J���K�������e��a��	8J!s���n����H�4���q���N��֑Y���y ����W�z	��n�W�l�������L���|GFU��{(�:P�I�]I�+z���c9�^�;h����|k*fx���6��r�0��Qb���B�;s>��������t��C�lE�P����UIZʣ^����#G���C�g��e���:��vb��a&��7�o�"�G�,,c��;���T0OZ������G[���۸�x�}Ӡ��g'TCD#D8�����9�l��/7�+�,'൚�Cy�r}xpi|e+I�_���MC��v�X<3cH*�;XA^̎�j���gr��D����s��L�鄗��D���k���C��~�97�qbN�W?DĒS67��5�w� ��0�uy!4T�/��b���� ����'kw"ˮw�����g�KF�.�E:áԹ�|��R����y0�T�ώ��4{y܁��zk�8<��󚸑�;"�}�a��U7ΜDLmD�]֟� b6�"'�W�+i�t���:��V�w��V���f��q�S���׺�O�"��6��;���:go�,���V�+��t#��~*����?���\�<n*MkE�	�{�k��d����vޗ׫���˵���q�@�W~Hu��1��)�hrR��VV �:3�e���Z�j�lvŧ�s��#�%o���U��}���S����+�N���Kt�)�?z�0��?�M��v�j���_���y~$����o�߂�}W�~�Q���N强�� �cy!��u�"m6�:�ԟ������`�4*2mD��3+��lo�qa�f��~��(�[��/k{��|a�R��y�c��"�
�rCw밫��Rh�d-�Ѧ����ve�h���~sb�l6�/�#,foÓ���<x���36��+��V��l���ҦbY�*�Z�>�R��!~MC����g�ԙ�uC5;V5h���𨿛���4u�ӽĄxLC?��4����g���c�rn��5����ݬ�]�7Ý!.��(J���T�vD�#�8�2�ݢW�,W�H!�|X��]�x?I).��������m����ڞ����J\�@;�_cT_��C��F��k��T�Bi��_	��wMX?�h�9��݁0)@��{�<vj?k�!|�4�IM��!�hȏ$�tB'�u�+X;
�(ӽ�����]��ܷ;!�2�l���6B�MO�L�P�ʬ�}�V9��g��r~:�S��PN��z��9m$�L��u���W��"V�D�w�:�����T���
�Bk/�L�ґ�ty�=�D�rBa�'��N��Z�j����J�C�d�?jH֜e{8Rv/�'V�U�A
�O{F��e�;Ĕyx>>x@!��ʁ��|Q�hO�� $F䟓
��]�t���IE�f�:�F���hr*�,qʑ{)O~�9�#O"z	X��Z��*�`݋Ta7�z+�͗��g{��җ�؋��КV!-��ҁp's��|���������C%Ae��wA�=�Bo:�z�Ɲ�}��K���b��^T�4���ٻzں��w�P6V���\��]�ñx)���;<blȵ><��<I�J���5-9;F��BC��o��:��7�uD�ۃ��x�D�5[�}�O�8�͗�E:v���\����a��3H;�|�rwU����-����C��M�Q�tKa���XM"��I���1�Wk�$Cۗ;��v�w56H˛yjۇn�}s8�Ϗ0����v����fw��z�N�zh�� 	X��x�M����*�̓�+T���(\c9w4�u/���dˏ0�P��'��p໌-���Fo�"���J��ց�s�A�s��}� ��-{��� b?���|�m "�1�A�}���U[ ��@�J�s�t���@�����3�Ƣ�D�B���r�2��l�P�"����6�2�p�'(�� -�rYK��r�y�ԑ&��j*ܕ6�Wo�]��6�@�����"c����óEp���>ވ��_�����9�X�4?�äg�GAA졁��&��jQ?$��1�D����ו�9�]؇�WN�I0�{{,d�ؘ�/�x���V���ը��7w?`Q|�@�m<�p�,�nOX�%�s=��b�"�aY����B�KO\%q ��oqU>��+����d���X������Z�v�H`�-��):�3����,Z�Er�r�$);]Rn���4��3�������u�tF�uwJ+�i�q�mD�jܯ��_�����NQ��&.C��h����p���O��%����˵��U�E2���VOs������}���N�2d3�����A����/|�.��y����N|;�+�ȳ�Z��!R���/��E����JaN����x�fg&��cK����ܛ<��.��tƪ=ļ������S�M�b��Qs>X�|��T�`a�_��k���7�����1X�����{)�1����h0#���f#�����]>���L��Ͳ��(����^w���7Oy�~�Fd�i����x/-� 6�8e``R�#<��-{ܡC}j����E8�  QX�+% u4��徵��� Ş��Fy�ss���8��q�����^YO d�Ӂ6WQ�xP�.�]~A�v��N;.
��~�m�y�iک|�v�rE�L$�Uv8B.�� Jn*�c�g��V��<�	o���%כ��wOȏbh�ǹ�F.jc�ݻ���;V��g�;�������]�_�J����GF���c�g[H��D��M��";I:1]7Mu�L�s� $bFZv[�����+`��d(������;-�S�"��@�I�QƖG�#ʋ1J�`!�T��Ґ�˒�-�˓@u���$��L���7�E��iU�f������*=�e޽_���Ȼ�\��@!���I6b�2���f5�8G�� 'I�p�1i��C�%Ռ��s�������v"��,և�D?�D�R��;��a�$��@��� 8�/���T�c'9w
����p1K(��j�ʅC�"�M�j��o��i����s���m%A���1�Q)��9��$���L]��dX��3)�������4t�BO?���[M��я�����S��m�;c��!-�MH\S�&��`�φ1���7���jh�o���Y�˹����G��<����^W$�AQ������S-zF���.�w�ԖG�a������,Lc�4��S2��gF3��WyT��J9��;���&T�6���� �c�`��;�03��k�����ړ��*��a�7�s�Į�|�wc��J�t}������ʈL�x5z1�_I�v�������SI�1+�o9�Jb�;*�l��T�9j�Z\wr�$9��v��u&��գ�t9�K	�;�; �c��`.�H���:L|� ��`:�Z��<���7hhRc��\�5�^�
���(Y����X�d ��>�����(|U�RD���ɬ\��)�ޗ���z�b��X��1C�p�B��x��ĭk(��<�����<63$��_��D2zTy
J]�[��^�)���ZUؖM�x1���#=�H	J��9�XD6���f͓!�s�m�#����a�G)�����14����o2��-{�i�acVc��}��	��X��Ea�a
��&�XNR=#S�o�[>�*��amxg��//���^>8D��~5µ.G��1u���t�����j�hj��#���M�X�[꛱HFnn0g���P�:�a��0��7z���X!݁-?��%���'ȷ�|,p�+��lhz��8�+̥���oP7�=[���+_F�2����8l��l4�Ud�ٓ��~�-�1������aq4oq�!oEm���_���I�(�/1��⨛�0�	�G�7���Dv4N��YL(�v�9��4!_�� ������`y4�/%c���r͇hR
��pDT찪)��k�e����4���>M�#��`v���0fh�Z�&��l�)�0��qp2A��X�#��u�k:/��Ze�Sa�9��;�m��������~�>�杋����p�$(HsX=Ey�����%�@C�
b���̖_[�B[7����'>(}0J�t���l���0̄�"�й�6D䩔m�F�j4Β��HvuZ������I+�4�7�^]��A�'##5�7O�M�T]_�d3��6����#8�h�Lou�NE(O��Ɨ�0M���3W�S�,��C#=C}5�ȇg�8��R��9�rC?���KE�V���2����w.�>3�g���#�X�E~jnJ��r�|��.e����b��n��_4�<Y%��۵���\a:�e����؎��_�M�Ϟ#��o,���G�z�(�� r���	��
������?���
,���@VZX~[����T��=�;�kl5^A����.�0����vR���z��:���,�Hx����']̜�oyK/e6�	Ke(�:҃#�i�ҲZr&�d52Y�7%����[ǽ�N��_�-H���!OH�����x����C=4
^�\��UN��q\Q�9�9�iJqG
�M�_s�=�>�^���_�z(n���d=\�0���1�Q8�쀢�f�A(�aLU��,L���<H��ۖ@�+��P��J��� >��BAr�VhL���Q$BCk��c���XD���yA}�î���oݥ����i 1	�����`p��/W�LH�a�vϟ`�}UoS�4N�-�å�>���W�ݴ���H�B�=���"�Zr��G���y�&+��q����m�GylG=����%J,����fG�v����>�&O�_X�D̈́�eS��8]/���0�tSk4u^-`���&	�\G��Fہ:�b򨡘@�>8P����g��"4'��U4Q�AO�CR1���>I�|�_T�w����Km�*3��GI6�0\՗�Un�����ٔhՎi���y|?]ws�6K�|���k?.]�g��0rع	���'����z��osq��bl!��������_P��K�r���s�x�N�o�r�݂I��N�<l��S.�fΣ�܅�S�knWI��op���&�A��{ԁo����s��#=;%�:���C�<��6�h�b+}�Jz���
Kо�Z�V`��10���>�w����
;���$�s+�:����i|G&�W��V��D��}?-;!FW0m�|SC���Y|�Y�n���8"���f7��/'�^� ���ص�P�mnME�}P��XWK����\�ʄ�oj(EUc����m83��m��ah�m�������@�`(K��L�L���x{��e{�b�ך(|�p�N���͈ɧ�B��~ȴ7���oS�s��{œ�̳�$YO]5��Ŗ-�[�Z�q�d��;���(�}���|^�@��q�A���@w6�9����#Ux@� ������������g����Y۲�̸���:c�UM��²yy����(�~հ�����e�^����
���èp�KLqk�n��j��w+�1������c��˅v�S�Skm�B�)�Ђ�#qf��i�55�ѵ�����&Y���U&�z|�7g�4��H�#�!}}<.S��v�h]��Hǖ���Wb]]� ��p��I�g�F�n�Gž\�oT�!�+�g��܍"_�%����2��țF�_,�1Gr�<�}��xk�X�K���~�r(�d�	�{Y�ho��G|fN���Z)�Ǧ�#de9�\��	;>���f`S����EL��U?�S��B�7��e��p��~w������SU,C�_�]v���jw�!��D���m�9X��i�@H�WH��~�����m|ʍd�~s�#������כN��><"/ �m�'��D�$���\� �?G��̙es5;�b�~3���|}���Q�l~'o��|�����08*)�Y�%��@�߷9��{ŉ�%V��ƴ��4����i%��;�y�N/���:�8.^����Q���f8�� 4d9���I����.{��5����
\v�y�������,M@�=]��f���hy�ԦպF5�����;����uH����I���:bQQ�9N�����ß��|�Zo����հ��k��וu>���ǟ�h%d]ٌ��5��v�	�u�i`�oU���|8�,���v��|ђ��\�4�LUA ��1z�r���!�g�Q�I�6��I<]�����[�.�9ʪ[�����M�f�yÕ��q"�Q(2�F�	�����˻2���·���+��bv�|���X�o��a&����x��k,g��d,#�K21��A,���w�Y�J�l�PP������JHj��-f�q���0?�6i�'Q0���
�%e���Y��f�~��w�c���;�!e��3@l$�r��׊H�ټ;�x8��(��6����Q���Z�Sl��X���ؑ���;�����!��Tj��]c[���4�+�ޒ��d��b�Kz^�ļ�=^�#���qh��n�Cm��c�r�E3�<s^�9&^	R���UKo(�1�D	�����z�b�dI�$��j�����>��E��@�"�4س��r�X��5˺�N���3��b�����n�v�1#c�^x����r��
�T�����OP_>^Y���T?M�EAt��{F���֧(�~�+�� ��Lp�V�!
)�t��/[Yo������(G��8O�1��Vd�1���	4��! ��w�tz�t��cqB��5�aZ*�jU drBi8JZ*<�f�QԮ���;{0zSQ�1q_�%S6��ׂ!'����ȥ�P�q��۾֡���?E�i_��x�Y3����e��u�_.�>�(B��D�&�X�Aj/��$������TTĊ�|�EM�W����/	��,%�'Y�T��?�i%�P�}C-�y�8��[ֵNW�+d����٤�#Y,ꑭ>���2Fd2c��YݟF|����L:*.��b ��3 ��i!��S0�!��'y�Y�*!�ɑ$Pk����,�]��������|�T���? J��NH��E�5��E��.�>��Ɓ����l�a��Oh�a ��ȕ]�ќ��>M� J#}dÁ�T�00XE&@'��L�V�X ��P������X���d��:�O$�4��&�0@|����r����x'u�ǿc�dM�yZ6�z���fZ1�CI@�R��=I-T#*�$3>��
�9(a!��	uZr	�ʨ˱Fd!� <=DQL���c��>/�Ke<�)�X��-�_9�Mit�a�PkSjjLh�)r�K�uW��
F��R�[��9�G�ɝ_ğp�)(����\������Nw"�����Qfrg��7d�y��:�S�nt�� �=�V�<]���b��x��2�-�)��Zp^��J)�D��<�8UT����H�+�p�"JC>�Uy���A�,���b��PX�f�D���:�h��ݎ%�S���eG��jUQ�5KŎ�KV� ��gv3�K>T1E4g��ZF�磙~gME��h�$&n",����֤�7��ݙ����3�yz?��'���g�)�X ���r��ꆪ���*.���琐L5��kƪ-��:l�b/%�l���#Ʒ�P�N�[�*ʏ��@��Z���h�-�x�)7� �"2����V�L��/P�~+7���a����i��Ԇ@�����4��JE��N�.��g�|r^��g��î[i��'J�s�<�p�~��*2O�F���~aΜ�g�Θt��@����jrs��j���F����8�,"� �?���-�&p�"444 `�B���\W�]�dB�=L����*È˔Ýd��!	G���)�����G�;8G��[�Nl�۞L�L<�m��$۶mۚض1�3�w��'�ԩT��;��׷����^)z�d7�Zt�M��K�7$8���\B��������WF�%N�DS� �W��gˉG��k�fz׷�#"��dz�d�`X�������wM�ݑ8C���v�6R��-�=Z�w�jڻC˄��!q��@҅2����5�a,e��f	���G�z�oˍ@��"�����#���Ju�A}�9>..�ޞ��'Z8A�Z��tx���G��<��d:[�/u+�nԉ=����Jiee�d�8x���_��$�P���0�mb�!y�9A!�/�S�t�
���
�^$M�r�a��00 B|�k177���H
�%nh*L�v���T��dtl����RmtrS!@X�б!�;" ȑ�bM�(.-M�׸'	��K�L�K}�Av0�$��G"'���UW���LA%��eg�{�`G��-�����u��BW������?�Ч�4xRcLW��w�[|cD����B��y�� ���a �T���D�A11�_�Ӑ`� BHJ&����,T�S����НVſGW�2����s�ϯ�0��:`�)��j���)��Z�Nz0(L0��7�熌."4���p?&�>�,���O�x@���O�C����as)I��7��Ȟ��`�K�qN],VM�!���N���DC۪ʈ��$(H{OJ|�+fۦ���o�����5����q�˙���W[wnM��It�Mny�r�U���AVS�"(�<+�ᜃ�t<�����]�xu��������锭���s�p�"nw�D@�nS��SL���i P�3��M%:p�\7TAE;��jR#���CRwx?-dp���Zz̏&0�4t��o�r6���}<O�j��
���7������}j�NM����'b �YDpz��eӝ�����#��I+���;Pv�'�e��󖢥�~���Dڵ��41M!+Ɋ�?���5�i>����J�@�1n�������s7�|A��O�A� �O�P�-�k]%r_�ȿ�}@�<��k�p�>����rk&�ҹ��ܸ=:愶y��9�QL�-�,���s�(a�J�#뽆2ಀS(?႔��9�"Y�h!5���$��E����h�y��6���H$�(P���s�2��y���Xn���c:�y&F}�)kJ+�r����-})۾�O�,��2I�JbP�\]��(j'�pJ�̂������e�P���w΁���,rU׭�rx���M�,��AO��$�
�X����A������z�;���8c�g��-w6�(��f2�+��עc�3ݞ<;2�J��c�����)�K�ժ^�S����|m4�y��	�������/jZ�%A�bnU��	nJ����Rڽ׺����ng�O��/-���o�N�]	�'���Jܓ�^M"MD���	�ь[E�I���<v`�o��f3ny�9���3/���Sc�BfM���1N���4����ު͇��{��5<=�5ng�;0��{��/ 8O��v���?r���r}�����AwȦ �)�����`���=�ʛ���'̝1��J;�������:yH�ߙ��r�s���,��؛��ճ�$�σ  ��'�_D��G��@TQ'\�ϊj5�V�8����?��e$R�7^2n񻽵�U����[3RK[cI������կ�<�.��������5�7g*{ktj*?��h6��S�#_���9�� ˡ��;��D��~�"��JW�G�����KR�Q�z��+E:[d��E������,��)��tٰ��ӏΆ�d�~�8Tf)��uxh��I�k�q��4֩?N�c6��^\Y�u��]$)���K@5d)m�X�C+#4�R��[`�T�����0���H��g�S�!����r�ѶORc�U�ժfG�RLm�����uآy��T���BqdP� 4b	Ԧ_1A�:��$9�燀��L�y�;o��[o�Ȱ_��r�a�^9	���NKq�&�0��$��NmT�����5=�����M��y��X���r�saJ�
k5yM%���d!��5���`�8Z�.3��ǄS���H�P��c1��݌H ��nM���0�ڽ_.����[��W VȞ5�?ʜ���/�#zp��"Ew��&�cE���'�PI��4����?6�n��
��a	�"Ǹ(���="���H�{-�C���B����)�YO�j�-��7$�B#�(Q,8HF8�D�F8�`��R��	υ� �#3���:�q5�$�j�ҽ��a��tx�n��{�<^���QJ�@kw�'X����p@�P�3=2Q�O(Ø�0$p����������Z.�6M;��k��o���#; ä�C�^�ls;K%d����x��l�y�-�Fu�
�寴-�T/k{G�U��«̅n�z��-��m���L&!�Hǭ!'(U��)bte�#��H`�g�	ոi�����N/��(H��grњ�A��X��"�B�� ry=j�I�互�}ۢ�?@k��u	QBw�[i�z�;?UDA��N��N�l�{~�9�k������:>Z�6��I��
���`p,��N�ǻ�+����rWv�1��O��(�������3Ո_�u�I0+M��~�+B������~�R�y=� a5<*t<��D#*�S���N�;�4^�����D���&'�3��rN'�B�m�@�v-��rPz���0�(r(w�Ǿ�E*��W���3&~�Ab�[i��V���ѿd�m��a�b�I�a�J�.�Pi�^������m� ��s�t6WC:�3�!�m^G��lx���.�J�[WO���0�ѥT`(�d�#�q�q|���R�� ﻞӾ�{B��z��f�q�yY�M'6'�«~!7�&��ϔ�tCȒm���k�E��ԕ��#�0Ps�W���bbx>�V=��=�n=����&Uz}���5�=tc壼�wC~}��Q�ߤ~7���>�4ːW�7W ��E� *������q6��)A��A*���]�RV��~�JA�C'�9ߞ���rșW��U;��*T�cԀ�b���Gĝǐ�����:�fWo�N�HK-y���MMd�q*�忞>���1����w�pq�[%̞���#�_�����2ZX�>\
�w�J�3O�����)F�ۡ�UT3���<��Rf����"p��RT�0�+Lǭ�3����od�P�i��Jwp��"ֻ�@��N79�ņ,e����~��)J������v�xY:�&�-AFP|��F0gR4��$�ȓP��?YL鸪��h��8���e-��7�h씵\&�j�:k�*>��l�T����C\���B#�F�!6ϩ0Jh>N3��6� �H��nO[��6Cڶ8�F�JL[>���;ο�h+�0D�g��`�����@^�3�͞s��**���_�h��=ϡ ��4M}�� �s���a��LE���DNZy/�A��+~t^*f�ʇ4��T��.�OˎY�������,��(�E�g[C���4i�hl.�M����5O�����I��8��PJEwx=�gz�k�@�UF}T��Y�Ш(�� ��r�U�bJ//~:M�^�*Uؓ>���r��FZD�}K����9wmT2RnK�Ȝǯ� �_�l����ƣ���/2.��!����
y�2�V\�m�	[�'{�� �v�*Zl�?�����oq�K�|S)YY�ۣ뛛�Ώg��؉"N�)\5�)���b��]��~�{��?6��\RbC����
2ѯܰr�������ch�U�b�+u��8>�ө�� ��e��y�7�k%���s���)
&�@gp�ٮf~ُ��׍��xf?�<���.$���O\���b���ܑ�����)����{�T���yhS���yݢ��[O�S�5"�<y����딁ɜ�.#��Va����֪��
f�`}\���#���	L_�hEhŵOZ:T�7n�'�F�]��S��ElO�B. ��JO8����8Ӻ��z�a�����Ew̓v��ِ��*�z���~Ҥ�޲!Ve(����q����.=2&���\�E)C��j~A�Wւ_u����N��g�W:|	Gr���%\�j�x��s>s��`H�����<Ʈ�6�X��Kz.�	.S���&��KwҪ��kk��<��u�t�����HLy�����YN��]�d�+qԅ�-�G)Ygۓ����q�X[����G4�Ap1���w��B��O$f�9�-6Z��Q����S���1GV!>�!~w�POĦ�����������+�|mp�f��/�@��)�*�'�����$����Ĉj5�ua�q��/�,�Y�����\l��:�/ PU�j��E|c�bHK������&����㙞��T�D�j�)*��Z��^���gO#�t�7A؛:
�|��F|Ԁ�Ä��C��@)F�n>�ڄ����>����t!��Qw����TԖug�����X����A\�I"�w�tx��D��]V���
�4�1߲��7��h�5kt�o1�@��i��^�����K�\�u9qq�;}eFզ���*�b�6ł�I�i̢(�Cre�`H���pjۜ �@��qe��Q�`i^3�!�V$wS���V���{U�y�� �Zv�<�Y��"h& ض��\��|�{}ɼ3�%���avP���P3H0�Sj�A:�Y�Ȗ�{;ׄ�gO-tO��Nv �ݡ{����_� LϏ-\��XGX�N�"}��t��t�
j�X#�!7�a��o�5J�+���]�۰��:!{}��ۿ��k��vٷZ�-�����>��y��y��w|-�b&.Ī�8�٨�"	�H����b �l$,�G�
>��7ՍF��m���Ȱm�h�_]�_��Pud8h@�~��~T�7�e]�dltHQi��2Z� a�lU�1�<UV9Ȁ�^^�c��wB}/��,�~D�.�$�Za7sR^��uםJ'�cӾ��5`@�:��[�����[�6�x�����|P�& �[W8A=�e�	zz�jX�*~��HJ�
�ozȱQG	�G�X�Q����H��}#�ဖx�ʸ��Z�P�u"
,z\���y�>����mx��\��o6����z4#��ޓ�*a4M�s�xr#���Ø�{yu�"���CL�(��˫��LE�We���ؖ����39�֖�3u�s�YWo��g�j8���P?���׶|�M��c-9���Q��f��e>�?-�#����93�}LNJ���4tT"�����%��x;��M���;lh%t��%b��s���\���=���;2��Î�ﰣ��=�(�	��7���Ǫ�!:���Qs���YY�Es)W�毷���k�
D0��� N�����hk�ʇc��ks�>�� �Xy����`����]�؈�KƗ	����Z����==.�h��`�H M۫h3NK&�O�hOP�X�T�ގ����jM�׍U8_� zA,8Z8˷���}�RA��c���,�s�}�oi���W��-��e|��d�cmפ��]X�i�w
�.�M������e���I�:r�=nx0�w��[���aA"�|_2���v���;Q��O1 MЈYp�?��zA�"T�/�Dbx0��F$**�"V#�D�=LI�I�3N�XC	��@D	yE&�����#�πC��[iy��L;QG��)a��F �v՗�(@�XV�0JI�)�uM ��FB� �E������lЪ����`X�ӗPJ�D[?(o�;:�3L�7���9�O�0
�]C�1���Ֆ=}�	��ӫ��^��R�{��L�t�؂�)�E��k�iH� Y�Ux�
F3$j��u9@Rk2���ޓ��G�%���,)�Ë�S����,���Kie�8��v��Ap�)X���f��d�0��@����N>	�<]?�``��B�ŉᴣ��ܓ{�2K^��m������q��謝B�����L܈�ⶆa�P��߁xo�n^��6��<^���K|���}�݁W?���3�:�TH"8߆h�J�Wy�Tw��[\�?�e��@�w�%]�Tdq��'�QG��i*��ǔ��A�8�QDR���C�n�n�@Cdy�vݸ�%$$�g�\�ʛ�P���<=3�	D<(e���/9���<�(V��}�D2����L��rL���������(��S��2�GX��p2�b�셇�E7�/r��c�Y�f��GI��!L[��o�k�)r��z>�:�/4Y�wuc1��mp(4g�"��W��r.�P��/�M�l�2D��ֿ��EE~�A�+Lc���7��4{��[j����U��84���17�������y���l�l+ڟ`�����
����)"��,���O'��ε�PRo�]��@/W���թ�����?�vq�����sf2�琣�ۄ�v ��@����,�~Y{)���)��C����g6�J�qY�	P�Ы���r����lo�2�ϛ��,Qt�tA{�6����`���彤|@���|��ha���!�AK��h:x��$��$�!q�G����U˙��Մ��2�	�3��f3�K�z`�#;P���dmփ��qڗ�f�����aQ]���c�:���S�k]^�졟��M��P����D�[�B
��b��VY?����a..��-���ׇl�A?�A����0l�A<��2�t�6�}v���3-M�-O�H���.H�ޏ��ʫ��L�'�`B����	�$H�/k�|�k��`�XdJ�VKgL׍
85�����"�Qp����n!zkVV
��j��PО��k/��غ�ۺ�oۺ�2��1&벦������AA�� #<�\�
�b���!� �Q^��yP�f�g�_� �lE6����5�N" �3�o`�E˯"�/§s[?�8�)O��2Dã;ER�Y���R�'��Ƕ��N�R4����Eט8�1�k�3T�'����=���ꀈ���ZZb�kRAX�V���~%���$Mml����`l^lDA��Ht��!���	��͎�0��a�_����+���L=�-m�*��pÙwE�������0>v"����-�U=� ���j�5�ga!�s��)�($�u�z�i��0�����ˡ>=�*}k,��:0��V��d�H?,ʳ�MZ��� ��Y�pUm��:27+V{��w�����.����@/��~�Z�@%�Aѻ KRc�cW�w�ͬh�:�l�Ze(���+x�E�<�&M�8Ɔ���gp�7��y���� �ث���i���3�?׀Wؚ^q�9<y�<M���,�k?���te�7i(�AԲ퀛D){fs�_!��t�+��W���g5��
�=� ocQ!��N�~E�8my:k�Q<>�8������^]�[U��HI��v�ޣ=!c��	k�*-��^���<�:-�KDhg��G�L�|X��R�YB�x��2�#1�L.��E�Oa:�]� B*ߪ���]���h1���U�S� �t�5�`©�:���mEl ��ɫ00{�J�Ʀ��8�)G½k�(y�?����lgr٢�j ��w6;��{�4�L����!iŦ�h��EB@e��x�粷�c�5����5�xY�ph���~�awN�Vy���F���6�H#s�)�!-��(�cւ�O&�eۃ�e�B󭨉�4n#%UUO��`��E�ā�3�u@ �1��p4�U��^S�!ihp���r��;������cҼ���/{v��$]�:�H5��p������Zt�&$힤u�φ�`k�����%��+g��)��v�-R^P�*�����K���;�g�F���<��h�v���[���f�|P�M$�Q����|��@(�0����6�m�>���{�q7��И8Q�Y
.�o���R ��h�Bĵ���st��|�Qb��?��ߘ�{�.hX�=�����(.���::��k�s����[�fE1z���^>�v9=��RQ��/���8g�|��t
���b��@�x�n�����9w�]LY��^�5�iw���*��,���m���q-�RVȖN�W
��3��C�<�/`f\�-C)��qwy�B��Seg��)��q&��Pd���3�S�Em^˚Z��a��8ˌT+z�ĵ�
�h�웠�fod�}�e%�MC��zXմ�����3���֢v#�x^��D�L'�ܼL�-M�n��e{��`he�d���W��'}�����)���V�廤�p-�cy�AZ�*�@�ig���r��y���ǟx�2p���zjq{�/B_�`^�G��!�����AF��a�+�VM����lbx{KRl;���K1+��.�8��6L2��o))ю!���z���Ao>;��\L�X.v�nF=`��"a��X�E���������]xї[ލ8��_sB�K�������Y��̵��U}����D�ƞq0oU���T*�,T��h���,K�z��0�Fw�x��򸾑�qލ2�G�G#��Z�u�r��M�Q�"ybuT[D���x}��5)��I��,vt`�s����'�}��H!�~�&�AƔ���,a`�r��k�1��O��4��.����i�E"]<`������ke�#�X����iZ�����ܠC�\�=j�g��g��.���{�JO�c%��~��%`hԾ7aL���ep�����y7(�
��`'�m�`g��=YF҃Z4(C!�+�g�����/���NC_�d�Y�X<q0��ԵY{����%�h�H�qɿ�K��d7������ś�x>�_p����6�%�qy��=��RQ���Л0�|%�������ƛ�}�/�-;�	E��P}���3ѕ�������u],�>���?GV��_�?�Q���B����n�\�z�%�Z{Z�=��v��^���;���"�W=�&p�\csR'Uy�װy��y[�<7�=tJ#�t���ɍ8��Yq�K�D�(:7�~g��JD��fپ'�,V��|qdG{���[y;Vc��Ʃ��}����U@�76=ӟ�g�#V!�dw�y�����D��kI`le8�u!a����������GZ��R��-��N�՛���"u3<3{�<��QT�Ѭ�.��0
��I^�K%����K+�I��O��� a}��U�1�-�G��E�l1'AW�ʪD8�<�όe�Z��i��,k%��5��=�&���cCќ3���Y�m����ug1�Kw�ԓ\n����#����m�ࡧߔ�A�� fo?	�o�`��>�-ZHru��D��ޫ��J]o�B�T�80|N5�?�	�7��Ej��|�-����&X�a�>�>��ML�@8�,���]�I��ke��K�ȡ�����Au5�4�U1}�Z�z�#;zpB;� ���0�����Kt35�l�����^͚��D�>w�
���3���v͹NсQ	��wF�P#�w)	�?=���o�%x��z����:oYh��6�֛�c
qE5��U�`���2��y��`s��}�E9�~' ]oo�
�֒o��/O����RrʛI|�tXRBҁ���Å	�vhx~L)��[���߾�G:{,�]�.$_�$5xk꜏�q�N���*b�3��I�O�j����R~W��N�E_����@��c�^�ZFϲmS:��5�*�2|.��W�@pL͂q�H�_ݞ�X�"՚����g�1��Yį��F�����ґ⤎X"�;ԗB9Nq��T:��ј�5�r6�J� ��mW�VΝ��V_~���a1� j�
�� Ӟ�G���D��d���<L��'��F^�K	�;s�a�%�  %�vc;�{y
A��a�,�-�K�tZ~bQ�H�"s]yu�Ԫ筂&7��ɻ
ѽ����"�/�f&P:T����]�I-�.��y�P"���t���B\n���#0Y�F3��Ct�϶�AD�{dM���"h&��48�Q�q��s�,b �3OOI_�NK�m�·T����z����mw�2c���	�;�%���s�9�Z $4�+Xg��D94�9�RM4(�Л_��?��3U~�x���J�밅����eb�4�dʀ����;�	�yD����U��(#7��[�(��f؛���
N���9�ԁz�?k��Eބ0U��]H12\�⣔��vf��X���K)�.:͏�7�ka_ӊ#>'G�a�Iǭ`�|n0y;oH��j��"��㎯��v,a���]��N�mc�}� �#W�.���
P���S*��ùD��ũ����rdQx�^�_)s�@��9��:�?�*y9���,�Y'囡��ņL+�ni��k?���O0��9�y�?�^�@q�b&9��4z|ϻ�GW|X����h�^_��7���r�k. �TJ����ke�af�y�̊���ti�,&1���<��Ac�����5��v��o�N�v�WkQ���u�m����*-�ɬUD�˝��`��款C����Q���[.�������rh�Lt�-��w�� 9��dTR�!��%A+�Cڗ]Vْ�B$�fށ��M��)�V+�ua���{��5>N#�Bqee�&��ZH��~Źa�П@��[���
�3�.��xe��;����wwo��)D����8B���{Z��N?:3�h�x3��pn�rC{�TZ
��Fy̍��RD�ϱ�6^�����
hX���P_�,V؝��'���Ʀ�����j$�3;�q���]bȊy]d�\Y��+���n��hq������-�E��c�Bͧd��飼�H�Ƅ&zo�� To��"�g�L,��X�)�Բ
h�gn`H�y��<����GR@։0���+�"î"��P��I
�X��܋�=��0����9%z���y�m���k5Н?�23RG�V`�9,�?�L2/U\����49`f+��ׂ[����tQm��:�J1�9⵪o�S��߲�:���b�AT���ɟ�%w;94�K�"�?EM��q�����4�����6tmx�Mt������2= `�� P�jX^ڈZ* 3k���TDd 5Ԯ��t�S��'v	�ei�|���������VNQ�n@�n���^��=���զ�Ǎ5o��ea�&G��!s���J|����{��)�F�8 (��,�/�?eWhl��ZE8/�v����I�r�}%]o>#((\�*#˪V&{\z��T���%N��Ö���ڱXp� kW|jI�\�0T!���R]���t3`��		C�y�����K�2�A���%7�[��	��ӫ6���;�&Ƴ�& �="(PZ+���\�-���5;nZl�#� ���ٯ2�:��A\9`��5�<�Rjꬻ'�Z+�o�������S>~�K�Pkפ�K���/���q���tހXk� +t�����BSE%�r�[�嵺�S��\��C|�K<�Q��E6�lGT���4N@�SJF.�?�5��<��|j�W#Б��sd�x��r7�)�To	�h��+�'U����ipf�oң:@k.�<��[���F�˙'g��J��{ ��a�\8)/��j�l���-��Kd44�]�	~�e}���gKf��.> >D�t��Wv-;�	�y����B��8����U{#6]����/"}\�f�}��hR��(�̚�w0ye�\�^K�o��-Nk�z�P��F��K'΅��dJ���|@`���V`�&[�
Rw7s��7r��vP��dĺ�Kwa�V��� F:[N���5(��2r��;���fhAa��#�~De�n�?���;
����fU��;@��>I��9�3c"?u��{J�w3rV��+m��)F�i�\�U�@`��MZ�$�l��2X[�-��E�V���⡁/q�ki2 �1�����P_<z\%��<[����
����v��!�h�t�ܐd���S܎`�$Svtkqp�L���e����&�4�1�|ֈ-�v3�db�71;����\ǒHp�zw�3(8�$��Аa���c�B_�w�A�$(���,��׶�hf���})r8�3���f�hu}�~�G7� �7[&^�04�ÆLZP�鄗�[+�Q�G��]?��"�}��u�0L���9�c�{gc�>���3�?�)0�(1u3�� �wsm�7��Z�wb()UA��VNsΈ]��tq�_�g(��j��{x��t�!�WY8�.��G;�����z��|9vo?�p��Fv88ӴFq(��oNNl�*^]��"��޿��nv��"��E��SSm5|"��ĦvT=bv�<���L�i��!1�E����(��]���r�nno�,�Q���g=|�fϧ�؏�U�5�\��0|A׷���YY� ���xVZ�!�@3��;� e�3�ص���Ъc��z�#gi|?O�x��^)�%!6�gO�G�"�n��V�gX��
u�.�v)W�7O�-}�΁ZA?9V����J��rfΩ���B�wqU�?n��F�5jp�it�"y
�fO|�m�R
�Խ�=��������8�Sӕ�0|�er��ዋ��H�u�iJ�X�I���5L-��c�d`�3�2e��^^S�2#�c #n)��"�|�xu��gz{;1�uZ��X��ҭ<_\���)g�D�����@��ո_�)>TA�|��`��L�i+��o�҅����8Xgc�K0��B���컷M�����]��Z��7��Ƙ/�����2$�{B>���ϔ�Бx��/�"���3r��?*�_��Z��e�Eř��� �G����*[�'T������_h�A=�h����������3s
�7�Ӷ�� �\�!4_F��J 	&(6)���K�Ǐ��ْ�Q(F�5᭼�si���g����c����۸�+�'ʗ��^�NpAs�Y�:��Z#E�2m`g3���z��	���P��dMbWCIP�2��Sd�HB���rFnlh�N��]'_��w�טh� ���ݸ�D�B�=�P����\D�E.���`q�2�跴��M�AM�Tp���5�������%�ʪ��C٥#br椊UB� ��a�7/��y9ό�c�zp@Pm�b�/���oT@�ș��55tj[e����%q1V�&�՜���(�����k�rl��}�VٟaAQY>���` �4щʹ��Qr�?���Q\N[¾�(V�� ��,:�o#.�-}bǦ,��,����w-�X��@�t|�E�Y+����]ʬ6�n�w�`={
���R� !��8�'{�����U2\�Bcf��x����������#Q�N �i'�?���ܪT$�	cM��#��h�7f��$8H�B6���\�.������ɒ׽iD���ϯ��Ӊ荃�V��@6d'��v*&��,%��6�9�U%3��*�J5��eȚ�x��[�z�gz;��(��#ܥP�b��C����7��?���q5o(ʹ_����-�V�_X�Q�p�}J������v@�?x����{|���˷wE�S���3S��b�U9�̓Y�P�^Ʀ�&�
�s��n��P�Ow�~1��g2��Z9����,��M�X؞ϚSz�<�Gu%��z��!OMG%r�O*�����;���tߤ����չ���Pu,�����nݡ��r���̈�����2�p(� hP�o��Z�6��r���\bcB���_W�g<��N�3w�ji���{t����Qt��GEv��aVI��1����v�6#�����Y��>�9����ڏP�?��z~{{���������3��������I��@?KL�kǸ3hlrÍe7���ԽM��N��ZY�f��(��l�x�5����.���y%1�G�n�H��J�����
M	��ʛ��&=������
+�+�����.ȓWEjtO��!;jo�i�VO�osC��ʺ�M�\w�?�^6�`Jw�q��J���!z�K>��w6C�XS�HG���ٰ��)�A�XJ�3g�`�������1)w��˒G���ʔ�6��Ė�G�]Q�k"�7,-��o!� p�v��Y�:z�Ae��𩈪��1�/��<��5>Pp�o����!��Υ$A	�L�)j�E[M�1�_\�덌��<�����=eZ�����qB�~^�;O�g���Uwp!J�o��&�k-�#.����r;���ɈtcK��lG�8Xq���5M�YK-���q��̙G�p<A�	��0�{ ��uEZ�/bŗ����*Mͤ22;�w	����k�S K�o�[� M#��� �B�W`f$�z�Q^݅�;95T|��:ŘX��i fZV�n���Ag<���PAiA�]=&��Ɵ�6M�n����Iz��7
RR���O5�ׇ[��$s1����k|����X��_s>FQl�{V9�o$��R�sW#�-Ʋec=��2:�1NT����RD���Ԙ��ٙ\UT1���&P5kX��b+W9��b/�-X9���!}�~}&�
���zMi�8���`����Ф��X\LS��eѸ~���n:�>eT�@� OQZ�
���@0s�?���[�A�괗QS���&~�nD��/��L>[�(��
��1�M|�6FVyA���ݔ��w��X�IO����Ӕ�l�Ϛ}��!����Z	�]�{3,�D �E�c;cn"��&�j���sa���`���?k�q�������@�y�Eg���F����Ќ�Ys��r��efm�h�̭t���<7�6������۔dQ�?:�]VP�W���B�i?������(�>-�p�p=#$�.��ry����j[W�Ī@�C���;>��t��/�(YNz�x���#����Q慄ւ�����\��	�֜��|ǣ�H
B��ɶ���8�O�6b�x�v�f�8���ŧ(3����T�1t��ߠ�fx�Jh�Z���%zc��m6Ӯ�R�C�c�tB��Jz|����������ٝ*7;>��S�īQ^t�Z���oN���,uΗ(ޮ�-�W,��6/<
]����?8��1h�j�L���O׀����,��}@��d�to�5����3=�0���}��i���DUbI�<>b�݇%?��O�"@_����X�;���I/Sݠ�}]y��h�d�x	�ͅ5m;5�����yϱ`�1YV���������|}e�#ۺ��_�D�3�+�mI��zh��˝A�5��Y��o� ��l����7�K�j�������J�.s�5�pQo�DeR��Bc���%����ޟ�����$��U�EM������� w �|'��ʀ�����)Z��N�h�jdi�c��]��χ xZO������:�]��U��J�=5anΐA�ͩ�aB�j���r�s��G)&��D*��2P�C�B��w`�
�Ӯ�2Vk���̆�D}�|��=��Fׯ?��Ա���`8�L���������fs(����33rM2<z)L(S�o���׽���+�w�D�7�<�����CZ�s7Q���)�+%|{��v����mS��,{����O�U��̗���,�z:_H�ꡉty�C��I��OQI)Kh!�:�PU�ʾ hS��֛�n~��%��q���U>D��^����z:�Z ��;}Q�}a1�n��G}튇7D~H�5Xh���x�C�����9��w�v�����.�|�%cr�]�]����>�A>��fD��J�'p�2����O��(�Op���ւ������J-�|SY�zyq��ύ�:�Vx��Y�o����5����6�K����>��{5z'�`p)�L��L����r�u)���R}:��h28��&��'=NJ���ݯ%$��Ba�)�#Ӎ����r!풪%�����K�*������ o+�U�q�0``dw��r�T�lھ�%c��<�]�R9���t��� �G]�R��V�6�+�X�j�nՑ׍����]�њ1�.��͞�p�~oN��y;��>��>�l�GLw�����	'.�ӓF������E|.�kQY�5����d��	�M�ھ�t�c�j��Qi��C�p���J��wO}Ԗ�_j��}��)�_�X͞^MШ����\����./�V�;k{�¾h�g��HDȫ0A��]t��U�2sl"!2䘪�1���
��:N����8|��j.k���'����s�Vw#5?9��u�t|����D'�C�⑺u�h�A(�%�c ;8��1]dTm��hp��e����^���5����9�H�7�wSf�$����@QZZ_���
^v���VO���j�n�7X\r�I�3�݊�sz#���]��P���gc�"���\���n��8�g���?���Eo����J���zv2�:�$��8P�Qyo%������D�Yr��h�-�i�Im�N_��SG��)���'�:���Rhhr�ذ(( �[����	��d��&�7�8���cߩ9�����QH�Q\=��K���d��$pza����s6>����/K���	.���[G �#�c�I�h�%����$��b�3y�+�+�G���Ԃ��$a�r���?^NkeY98ۨ�ŏ�]v�lNLK�d�A��?\�PM�6��ww���Ip'��ݝ�Np����5���K�{���W�Vm�L�>�Ǧ��`�T������(}����b���l�]�N����֜Ϋa&8t�/�I����+ᶾds�����3��[����
��;�;���N���+�̈�R�F��+�jx!�x�o< ĕ�H.Pp� -a��q�>��ۖ`�[�n-ը�,�_�w������;�9sa}�YN���hYٴo�̙9cN����y�/����R 
�ΝT�h����%�m�5T��Ei/��^��<��U�����b������&��~�7�g*X��L�P>��K�I��h��"��z}���_of;<��oC�X�Ar4�9���`jr2�|?��t�P�����|Ůx�mߊhÑ _NF�����\�����z����z'YA2ޥ�u��G1͹�T��R$P���M2u�V��	:}(oc,�R٣�]��a�x�T�B�q�n
9͈@�g�$�ݢu��]��=�����ݚ����T�'WU?���� �ې���.�6���>i�s���4bɚ�z�7��v�U�T" � 3�k(G�Ӿ��&�kn#���Y
��P����h;�w��G�t��� �E�탚)S����?G<���}���e�|�U❗t�	bҎkG�&�U
��<d���`�V<Jb@�%x�k�J�ɼ����A^���;)NH��7ӹl�k��ز.<}
����{� ���Vt�t�ק��󉇟
����_
w7ԾU5ѝvy���H��Ǘ����p腼��N���3� �
�h�X/��tw�4ެڿ��dG4�$k7?��~^t8!�[�L��a�k��"F�����B*0R�,��)Ȑ��Q�u�a��袲PY�R��t�@V 1S��'�(�vZr�L�N��-�o�g�,"�	�e�j��B�ۊ��Sۂ~0@͜�`8�M���>�Ha��E�eTßCg��K�[SA ���'�h�|Z�>8�omwۚL7i&�o��li��mn�z�>L&v(1�ʚ@:�R%�)c����l3��X��rũ���Gk�P���>>�YĦ_��T�@_�F.j9`����^�r@%�Q`��.��ѵ!���+M��\n�c���c&�ˠ^�R�/�$�C�� ��`\�ޣ�{���'��{}�ϐ������\{6�@-���8��|����>�*��������F�5���Ve�h(6ٹ�ĐY�&�@L���8���⨆~�\���.���aC��n�W�B��|26���l�ޞD�����%|>#������ rK�@cGs�x]iN�T6���FA��ɭ��O������E�������dn�ZsjMxV0���]�,Ґ�&����NU_&7a�ݢ��!�&����/�?^.�l�.8}\v���ˠ���ͥ� m��9,�5�Y;�CƦL��|T�#�(�����a��ڈ9<��{�4��eR;�~�);ZT3�ׯb���� �G
�u�3�Ɔ=�u� �r���]�k:�S�y�`�Z2Z�f~�_ێ�h�W���z��,O�Ý��Ew���̳������h�ڿ&�(�eO��gk-*Y!1��ٖ�R*҇F򰴔N
��_'�Y~����K]PR�_�#k�u*K��
yS�?_�f� �2H�x��{9�,"�6��gn����za��Br�)
���M���)�boD�uT�$�T4i�W1DBdt��~if62Ipj�MqB�x	�ټT�\&q�U��4�u�$��..�싮sH���?�AĜ_~I��{�q����V��Y��:r��v3�N�ufÿƒ_?��83Ctns6��=���}��S#�^��,#)fMb6T2��g�euI��Vev1�B�9�Ɵ����%`&ʎ\�Z��-.��,�M�~|���2M%T�1#����3d���g���dc����������Qq�ֹ��pi&!�:�M�r7��1A虌 Ƶ�Ý�����,l�j-���	�P����ǜ��:�Z��͓�<`�"w7�4�_;4n\T��q�yJi�	a(�n�3u�Xn?o��~�M�۝�\!\��jԿWm����}1�Yyk�ܭF�y�E�����Y��r��˟�b�&��(�84�����ZC�ǚ���bӟ�\�`����:���I���M��(_���V/��l2KTT�W�5�@$�(�h�OY���Q�*��J_�C�����MI$`�NDQ�NF�(si�߁Ȱ��,�/�Z���(*2����h��P��°�
��*ۇ�5���C^������@��A����:��q� �!�N��XK�ۅ��	��c�M9 �i!���M=F�mР�a��������Ba�@	��}��p�<��Ŷ���Q
�e�/��� 5ġIa[�cM�\N��
�t �������(?(��Q�/�+��O���0i�'&n�`�bV�]� 6oG�g�oH���l� g���3BE�jq#ږ�����u1�+�1'�p�`���7/��dP:��t�tX?�Qw8�W>�7���K cW���2	�� �Yy�)�q<z�.^�aL�$�G��ԙ�W0R���!@��W�<64���4���(^�Tg�x8�W#���S� d���W"я :M�� �2͹�%��ۄ<tX�x�v�z6�5�� n��$��7�Ǻh57�`h�����v�j�A����q�q3��nY,� ��rc7�jU=A��-:�36y��9�j�Yxy�"q7��0��0��98�����DN���\n�׋��y^T��⁐��)�@�٣�h�����������'�Z�Mqi����P~�N���n��}�9�����@�b�|���rQ��/�fs�qa�ys��L�3F��P�b�[�%{��N�}����z�XY��;��E���{��q���&(��O��MV`FD�޶�{o�2l��xN����x�O�6<�uU��{�����e˟��Ou>'p��}�`9Jiy>=���Z����"!߸����#��D�⿝����m����h1>%�a�ޟ��6�$C;�ھ�� 7P
'8v0m</J�^�W�#'��K�å�X:��o-��Am�5 q1f@�����V���A���Ⅽf� W��'���53V�pX�j[�ǚ�y�H;��(� �!Iwk��4
��ԙ�`bB��}a�����6���]���κ��KM硜�%T��d��u
*k��`ط����Bt�Cy^GlYY�;ᯏ�/oG.O�g�G��N�2��@�'���CG��zn��u͏.ô�]R)�˦�����eca]Q�]�X?��Q��;oJ�.6� Tcr��V�/��t��YU	�Xe��jq��O�ᯞ��yY�0ga����������
�h7QA�Y�-%���!��.7�#�[�\���8�8^P��c۠T�8Ý��d*�T�����ݖ!��\��b�H��}�1^^��U?݆�ubr��`Z_����c��-�m�O�!
�Еￕ*cA�f��QKs'f�[y-�R��> ��Ç	2�U�5�c��~���b��|�)�G�L�����h���-X!�ƒ2n�0{��?$�s���z?'��i�XX]狂��6��e�]�:�.^7�f?lB�p6Z��6(��O�y�)�Ο��f�����p�Ѿ���{��A��Vd�VIvB�%/9i��;鮽t�p�GQ�L���/�)SR5[�������]��Q��S`���S&��뀫����b�5�%�"bMض�Q܁���E���ع��Q���id�!mr�ag}D���X���k��x���?�d�}%�>��"T7�r�A���N���χ�SUG�X~�q�T;�y8xrySD0u��ZG��6}]�=��P�ӳ�+�����;�Dux+	���l_��!
�3������.?W5=+�\�t�6q[��N�9���?�0���v���v?���j��h���j���j�߈�`�W�.stf�/y|�Aq*R�/�'G���9<v��Y��Fi�6�;��&"5;=Н=���_��wژ�	nV�`�'#�O'�VY��߮ZUA�ŌQy|�hu���Z�h�o2����j�N��4�� @��o���&e���'�����}x��b��ꞓ�LPw*^����L�):i���M����;]*�u�$��*3z�7.M�O�ȹS U8Y )2����)O��x�f�E�2+���k��ꔄ^]��ݡE���K�U�&��=� ~J���u���5c���^���ӂJ���6�	����I/<�;+]G�6�Wmq�ko �_s��/��E9���<6NZR'��@ax��ǟEK5Ê�y���dO.������~X�IZď�n��Q����r��;�v�M�{8��͜Ų��1/�K�p����$�痀UY�S��_XL�Ȓ49�zY0����6���F�P$����2��ƛ�QN��Y$/���^l'L�l����^Z�N���	�~
��|#���r!<[ja}|�NV.�ˊ�H��SD���MT�:e�0�O��4&W���]j�^zf>���c�˘������6�( �i�mp#3(��&�O����̈��l)�P����DK�b���
鱃��=��ND�tc>T$��j&{�f4��jB׶�!Kp�����>�Z��v�4sʛ�Zz~ځ:�Y�Q�}��`�|��%�0�9�5���ȷ�d�{Tp�괕j����d�P�.^5]z0#6a�;(xBw�#ͷ&\u"��ڡe�Y��Hg������44�	Z���*I�/�x��%N��傢�w�'����i��	�;�AT^s~�����h�F�Kp��ٸv������GX�%;i�
�ڵ��\ �����]�VP����+��e���l��ͺ�ł�b� �g�
�	m*h����e��sTG&r��-�F�Bĺ%�|5��w��P[�HEJ����ƻzwHU����K�x;�g!�Ì*��ݑ��N���|��h�׬�jB�ྃ���i��3�{q'���o6}��r�,��Q��[jj��*��M�%ԁ�E����� ���C�Ksر5��9Fӻ��He��ޓ��hu�k��bo�͛���|�щ7�.JK�d��N����8����f�H�.�f�B�[/����,Ka(�Bz¯�m5���8ۿY�n�"��&�j]3�k&�b���J�J�W�<Y�%eyI'�3o�$��e�L\�iD1$�}�y����tC>e����k�%:��؇ƴ���_�����ݘ��X>Ƴ��&����r����(��]�^��p����X*�y�.�Ω�q��W�����xE�����W�T"��?��BxT/����d^�x�b�% A	�����`�LA���ب��d��N�DE�\����`��0S�Qf�ƍ�cX��(|���G����U+s��u˾�\F���y7���3WE�]���0�d�gu�M.��J���F�}�J�>��(Y��?=�<��W�����j�ޅ��#�0l~�떜^uPTn��V�
�^��y����]D��o/1���;��Y|���/���I��(q��^��ZGp!/h=��ͬj+�~Z�B�TO�|y�c)Ops��p�%�:�M����%��;��ͫ�L�֔5d�L�������|,|�꩷Fc�!H��/\ډ�7C�̈ǜ��Y���ﱅr��'�ԯ��q�ycl-��?�~2��<���3P��;�whUµYĴ�]E����B�١mM�g+���Wu"�u)l��=Lee�yX9z��##sEY�Lӟ�-���~��54z�c0� z������Ji�����fi������jn��?��$PPz�6t�ĻUO��/����^����׮bMz���ܭ�N���U�fF���i,�.�$�Z��
<�F?�����o��-���}O��퀘嵭�����k�]���6��w��؉��+|^�QCe'M�S�>e2#vі;o��}'c�n�]5�����;1C���^����`�l	T����4mm�؆.mK{
��������I���� �}GHy��r���|9A���N�[
ݳ��8����K��2�e�ڄ�<P�.*�xb�W����Vr���S����]�|k>�r)��Ţ�r�x��.<?̍?��'�x�jƌ��e ����~��I��"�o�H�8.'���۶�����u���c�t�pү�ɐ*��S���;��l�}���lF�+���l�]A��۔�\����۩�_��QVD�������t�Xלs<�/��<�,����Y�~��>xT�����Q��_Oxm/M�����Z����&$����FF�0+�[Nz�7	T�Xv��(X��O�,�3��,=/i����T��xM򺡵XߙTd~-Y~��	��}����uR�
��p�����kl�9�U6�̌x^���-��{>X�Z��Wq4ѸЧ��u�jс���;�E������x��Mh��__
Kz'�,c��wrZ"�`�6�Ƴ7peZ�o�tdeȄ/hkJa�KT~�6�o���7�������ڻ����`�ɿ���J�9������ۅ��۔e1����9-���1���y}�1y-�5����e��e��4���I�C�@��yo�"��G�"��i��O����ҥ\4�ٿָpXN`>�@B/hH3D�.���}r;�5��	��aK��X�Y+ ��*���i1�ݗz�qĮz�8���Tp���n�,��'*�O(T�K\u�
D��%�H4�njuu�֔mU�,r�g۟��Y,��hO�;�B6M_^b�t�g!��;�P��-�z���$�.,>������x*�jzpsD2��T�C���Y:�y��@kUȒ���:��k˹���zd)��ok��t�yW
,.�v���|���ꌐ�����+m[À��*��I����"	�������ލ9�/.;�9R��JӔ�Y㣨�a`+MuyS?|2B�i�9|�K_���XLZe��F����~e�2X)�1mª�b��;����Vg�	]�S8	r�/St��,H��T�e"��-�56W�
��7/��o��[�$�U�(F}\�bL�B���
<B��K!��g���,���-i\� ��!�Jcq�T �w�Ŀ�?�!��\���CCi�Z�,�r�)S�<�����in��P�zw��|�}͈),O6����,�~y0��H������^*���� g
gƑO{2P-����<nЌ�ա������5 Uk���3;GFY$�����7�%!M�h�5�ܗ�5��{LT�*&��Lw�7�&pj�}�ͳ��?�x8�)����-�L����ū���8�j��a�=C�xT+���~� i83J1����)�ҳK� @|��M��I@	�fA��r����S5gHN��z����D��)���0�z
��Q�q*(�D?���~�lV�O��7O�=��K�v[�$����L~�Y�1@D35@}��'��7���? )j����fp��kh��a�Bu��`�<��Iv�����
^>����Kވ򌦗R��1Y�G�T����H�[��Q��~ڵ�d�"�Mh�S�>��cŦ�eE��S7�D��F��+��,�������bie*��?�-�;vw|3�@vO������_�=윲��@��,.=�q�oh���9%I��W�p��w�`�2?��,���^u��.�Bʕ?���n]S�����(�7�G%I��c(�[�Q1�Z��u{{�G�Ν�`[m)(��A̿�&'0��D�����A�+g3O (L����t�V{=����S�d�-,L�h�f���V^�0��V$8�=g�Bt�M�e����?���޳R������>�J�mF����q�Z��n��Q�P6
�<+�{d@ÑF������%�H[�PeW9�'#���]�%�3��c~��&-�S��6�s�A�}9;'�����kr���U����
�0��n71R&��U�TN8����A�ԁ��Y�e<�'��`*�SF��FC.�:e��<��<nd����D����yB��1U�d:�J	�BZ[]>M G��`�z��r�����K�������ҦoW�Ar�m�烱>7p�[��X}����R1��0D~kU
c�C��Y+�����l_M$�Yw4:֙�5��)�Z���A��21c(�`�V�I�5�K^�%�6|��P(S�q�}�-�h6UУ%/G��b6�o���B�z�WA�����&����x�|]�\:��C��Y���ڣ�v�R�B�}k �����:B9Q�C#�v�LnP97K
���ڐ'���	��H� �XL�i�ao��!��}z�,�GK�=��:��3�� �['T��I��
����i�ې���1���PDq'w�@t��1���	����O����Q_�
��%<8��1q͌a�g[�#ƀ�X��ԧ����tE.XCW2��/w2���d_�"E���|�EeNg� �D�ŽD\���]t�!�������]J��Э�j9��u�CK�]��|����
6J��}�m�$-��m�yM%uBT(��6Mtn{܃�XZw�7?���i��)�֎/wBx�p޺�0H-4I��b2�kOI��/�N*\��?���Ew�NB $�`�-Q-�����f��c'j��O�r�+�U�3sj��zT#�5٪�P��Ũ�Å��S��v���*_܎����AN�P3�����l�%ku�]=_;��$�
���z �A�Cn45�� �ǃ�|#*�����J@Ir�O�"��Z�Ѳ���dKC�I某�%�p/|�žJc�L|?u!�� 7�j�	B{Wx>S&g�ɟ��1��#{w�2�c2�-���(�Yy�_X��s����t�jL����0$(�0���5?^4x�M��J��j�})}=cH���kCdK$�-w"�	r�ñv�]j[Bb/�z��Vg̲���8�L�ispk�¦n�L�8)�����h���J ʅ�4��")H�eHX��l��m����L�e������Ӻ�s0��������7�\�B7��
F�C*hރ�����PCg�����]3(����ǉ��8��r2�ڕ�B��bV���6DT�/�=�+�V&NV��@���w��.� �C�Nn��Pִ�b���=L�sZv&����@����C���݉E��d�g?*����"z�K��xg�Î�%��T݅��Ϣ�~ ܎1�/��s�4��ٺ#n��\�G��W.���߱�"��e&'@�Y�Gf'F+�����0������(�gr9�T�Gm�;�{�fG.c�\�N�"j�nn�%!f�������2T3�!0�8��=���Ϛ#tbq58О9c,"5QqbA�S_4'D�M�{!���>�#�8Z�rWn6�<3�]��{��Gf�;|�b���'Fڷ��CB�%���Ɇ�5ﵵ�y��υ�De!n�J#�~��%P�D5��o�� ����g�,f��Qq�Z�t�_��d*���EX8��KhN���K=
\Ծ/s#��#ip^?�������B�G ��(���:xܕ`�:`:v�.��A.��_+S\�a)<�Q��Ԅ��\CG/�}�ق��9�Wf�)"L��� ܲ�X��/��*%TޝZq�߱
@�dq�?ŗm���#��@<�Z��k�kw�g�I(��4>[mݱ����%anY�r}V�V٧���K��@���U�����C��]
D3E��7��T���V���2GBԎ��[86�A�V���..�n�������x�S {-�DG,2��VM�| Mu&����*ȑ��H}�u�n���=&ꐂD�@��ba�K�M"�?a�S���P����0�v�)�w�l)	��a��)�0���u�����K����9�ޮ?|:��U}�x8��}N)���_����D��$��c�|�vzp/��j>��o�[*7R�*�5rT0ᴝ�.�?믔���3V�*����%8VUJ����f���9"�oz�s3m�j���� �{�����������	nI,G���98��fG ,��;�AgMP�=��U��<R'���!�Aȫ�SZv̩�ԔI���1`�l�~h-@s|��R�N�j �C
S�tW ��h�oD��D�=�m�����xz�gơF�"}�G�z��A�|6���R��ۺ�O �wEۘ��_�����i�n PL�&���R�^�=��?�*j~@"	0�UV�WB�6ħ}+����)�b_8�6�� \r���>��v����,y��%'n�W��z(kh@(��ť]�{�'��g��I��j<A		}����`�u�S��Mn3����s��&�E05MӰS#�F#�YLxdi�i�s�#�w�|z�0�&7�NPA�5Žߤ�����qy��k��}������2UtV�J���֣V�d�U6������˔������.���2�Ƕ#7�c��EO!ӛnlkty��k@`]�q�d2fF��(}����ʡWxu��O���EjyӃ�|
���R�P�%o'�Eܝ���}��{v��1a���}��P���(�W�Կ�۪�Ѝ�ܖsmM�q����$��V}�Z����c���Ыv��P���\(q�L�W��U;/Kq}�����vb��#���3ި�Y$A����+�U�򜣆�����P��7j+���Z`*?G]�;�V�!%�{p�ޭc�]AA1*�ڍ�op�՛��+����!7xD�<�w1޵�p��K��z�����.0
=�7&{H��n��IS��s���=/g۽r��8���������.vC�и#�	���+[�=��jqC��(�#3:�aB�B�����Vj&����6��^&QM�T�ϥ"b����Yg1T5T�Ŕ8XO�EP��m��b��r�)O	6��X!����A\Y�6�f�(��k�Y�a�oY��"�M�X~�Z!���}�w�	n�V'��� �r\��Z7����vzƴ)!��6��aN�L�N��zI~�����z��ٯ�ub���fDaBX��;C�@���-�f�^sbw�ۇS[,�ޚ!-%��5O$����,j�y��#Pn����#��0�K�$�Go]n�]gi�}o �*4�ܟ�I���S���c�88�]�4���L��	��?�|)B�q��*5Ǝ���b �JUR`���]]�7��[_Β��!�)��4��������w�s���*8���m�b9����������K��W��kl�ڞ��=�ia�X����tfkjB������u�����y2L��cߣ�uZ��'i�e҃�r���f�~K��a}��5(��H�����w�3���!�H#2?L�&T��rw�p�Q��LBB8PKݤ�L#��
�Bf}�Y���˷��A|1�4�mw��w�:ѷD�g��͑�.7�������Kn/Ab���a��)5J\P%8e��c�d닯@�.�2 �]���8g4n=N(J��\�]s$\|I�<��B����\J���"G0�ln։v18���s&�^��������ڄ� Ot9w"9n��苽���c�Oޚ���Cu� c�v�B8&B�0!ב9��~��^��_�q�Z9�ü�6HY�2Z�Z8��:,'м�q4�d������)z�"���W^��C��(������o_[��E3�uiב�k���A>B���v�R����i��Җ�װ}�6~���u�����:�OG8cwtQ��\�T={ʬ���>���D?����3Ӳ�:A/+�q���֭j�\���a�t�n�z
�L��Fi��O����kԃ����������AL�E������nO�ܑ=��ҕ���u݆`����,��yǝh�G���:P$H�T�,��hr	��>P1�j���тe(���F�x)��x-�N�{��~R� @K$�sR0�MJ�8�ǆ�@7e��c�"��LØ� �.�k����@��Y9�&%@����w����:��S������]Xkt�Xl��:"�<�<�z���}�vdd:��nl�Om��2�v�E����<����eGh�u)Ռ�����n����R�w-�w�%��RJ�䲥\�|���x�W_u���o�;W�4��� ˃� (���	��ghG��@�]P�����z�2�8=��xyW�?�R<95�[�+ڋ����_��s���q�}z4q� X	��5TP���������	�q���F��1����K�+	A�q������͛�0S��1C@���5^9�T#��ۇ$���!���3���s���8tn:�v�k����˴r"��ͧ���ϊy%;��,���ozB��D1n:K�L���N����b�q����-Y�EP�#��1w�=O��Of�u+)���n����ǎ8�=����_S��r����,�Ӳ.��:Oڝ�m���F�I,c�@�|�$4%I�����`U1���׻t��|�ھ+�̥=�@&<2��v�/:���| ����^�3����; ]ͪ��<�b����3���^�����xL�`d�r��c:�9Wg9ƥ��FQ��M�	NB��~+�����ig�;�-Sj&��^�x�}n2(���=;�(�v�%^o��X�$����S��=��7��@.ݜ��RL���m�jG+z ��i�Х�$\�B7����s�@���5�׌��|3��G����,���>R�^����ł�A�*gh;�S�iP>�KCy\3��q�Y �2��T�@��}�a_�!ۛ�t/��<�ܝ�:滄s
iLn5��-5��FP�v#�HN�I� �����Vxw��i�`��²<�'�+��m�EÚB�<9b�ऑ�c����`yW��"/���$�β�Z<v��.�mVX��A%!REk�n@2�Ab"A�#�<��2^�^[��d ���O������ڸQĶ�UΛ��	���p�ݼv��������0����B+���F9Ll�8L�6����#32��oU_A�
�w�1�m�04$��;�篞v�GP �'V|3rp�����^�*��16�_�!����5�%�t���+~",���pQ�g3�ytE�E�"'�\�Ѹ#�A��qю6dJ��K؜Y�-LTgꧣ��)j�Q�/㱣f��}�
�_�o�z��ۘG
�u�dĹ�β���bێ��wo�Ce+�O#�������>�͍�Y+Z@�nB��$yL�-�FM��|��D>@�F�O���bW�ڔ�g��)�.[�ZF�.��7nù
��|%�p��9�vz�>���V7ӵ$��t�������ɀ���ψ���2y7MY�!�((����'�曅 �����t�����y���eE� 9����*>�R�M.�-�B#Kа��i��d�y*�Đj�b$���
���|3aF��G�l8��@�{j��z&X*� ��[9��P��
��~/�/��<�� HL���W�9X����<P�P�������.q��G@�I�jr\���|���n��j��?��1�V'}�C
�C@�1=��06��
����W�v*e�;҂з��-pr�i�;�o5��ey}���-�>@T�k�p����
����V?�ّ����124A��ڣ7y�ە	��c` T	3&��!��G�#��p<���P�������M}Iq $���f�*�6C$-����O��`�OܜI�vyk��tc��+��ܸ�X�v�����+�ҒR}A���1,�8'����T��?(�~Z_K�j�����X	p;
k �>�ǕږlL��0�j;���Q[8����G�2������ S��NAVR�<�����
����y�7n�5c��+W4<��b�ٌ�=mK� ��0�ҴЂ��BR���_�T��>б�a�X��Qg�괔���Db�K�@<3l���6T����YQ�2	��g��ĥ��K
���v:�g:~����j�l5�>C5�ﳬ�����oij��Rl�l�i�p�y��L����^���}�L���d�Ӏ<7~��b�<Y���t�xT
��uC-�Y:y�QT�<�X�`��7/�L��d�?�GXL�|f	p���P��m���z�7�VfҸ�b�=���c���`_��xr��H�po�+l���i���ޚ���XH=�C�_t��D�cP����.�BMM�J�����aO���,3�+
��7YW�F0L4gn��;��
c
n-0*��xTC3	f���I�x �=m��\�|�� l&J���/v������֗������>�a��/���2��A���jВ��
~ �F�8��h~�C>8mu�a���t�Y~Q�q8nPq��A���	�G���A�hŊ91��;�����~(���:F[���^ۯ�A(*~��CЁ`3��3-����u�Et��kA���I:�C�wE@��m�vaiv��:gv<	�vFu���8k;�ݹF�u��c���GV�iJ��v��a�e��?��aM���0��ޛ���iV����
�zh�U���SUQ�5���b8�P���Ga�l��@菕��=�a�T]=��r���3awww��f�g���;�Ƣ����:������b�>3����g,n�hʆ<nԇ;ԉ�;����q���/	2�̰P9^���5�Y��A<� ���wA�,���6����/�74>O39�5��0$^|ߨ�y)>o���E���f�'��ۨ�bZ�h��C���{r��P�� ���b�yl��{�^�� >��7�ׅ�����f��qes�G%p��mGp �6v�TYY��M�������dw��|J�!')��|�zP[�����d��/)y�诣���DE�_F��R6~:����`���CU�m�Ŀx��.O�'��B���>J�]�]<�ĖO��J�	��f�kJ�E;�i�� 	�W��B/��D_�x�.Z�km7��۵��rVI���\U`�(�O���|�[��/6EV=�+��v��%���ܢ8`L�+�#BR�1zZ �"T�I~q��8!�5V��pi��38q��T�Z��Dr)���Q���s���܃�+m^\yt-×�lT�ч�3�|ot8ZR5�bn	2�%`��04�d�aB^4��{���U�T�Y�,�E�S�P?�/G�&��iq���j��	C$H�!*��s?P2Wr2vr�n3��C��SX���A�ik��F0�R�� ���)����G�Oh͑b�&��k��ς��E���Hg��H8
O��Y��a@��� ��j���C` �B��TJ�%��I���$�q�Oh�K
���?!��Nh�?�B�����{��܅d��Z��-
+#q �y�s�Phm���a)�`?��y�?��OB�lSޏ���s�&*}�5t�w��"��?�AS$�!���|�i������[D�jw����?6���UW�̟���k�L�`�����CR�[42h�h���Cⶅ?�R��2�5$��!3����ꚊH��G��(&�&��j�'f�)#K�-�&!���B��p�8P�~l�����~� u�"r��\�ȝ���z�B��7��JU	���5'�v�[ag��ߠ����
Q� �A�4�R�!'i�Qg�p�� Ɏԇz�N`i��Y�d�Kի�Iq'�P���M��Wq5�EC�P ����H�
�C/Ifx9�ǒ,V?@���=�?J-�\�>ް"�b�'� ���5�(���c=)zڪߢs�A�̜t�(XQ�4H�Ұ�����2��-� �=DtRf60K������#�}H
�M]i�/��|���߫�������n]iW�}�	_��t���,l��b�= c�+/L��0�!,K�� �� �H*��hPj����J_���s����M:�&ް�[0��A�x ů��6V�ǩ�7���Ö;�o/ w��/2��#�#��)����%W:��$5I1��(j�!���Q�@��$�u=��?���j����u����\l �o���l�+�
������T1�� ���ΰ���Z��[���_]�v���o�3��z���(*�@�L]%a7vR��*�;���7K;��}�ӹ��~)�R�c��[�W�WB�4[f�'��*QE�q�[�(wȮ���#�ז=�������v�7��TV�����:@�����(df��ޔ��Y{���๸~��p�z�y��+�avG�4�U���!��-����j�]��dg�>�B�Sbu�=>ڠ�>\��j1PY}���2u��;#u�쑞��<�:�x���q�:���l�Wj%R�{x[�^�ȃ�A�n�Dl�|��<��%O��\��u���6I���8$!��L�J�щ����u�_����o�}#<}}& )G�òT�H�q����ڞ��|2R�]�3�!��|����g����(Dc���!�	��q�ߗ�h���N�t�/�'�����EB�� �I�����&�T�5�(f���P��"�B4Ht��P�:25��ȅj�#�M�~�^��ܱ(��NC*��N-S5�&����;�m�������f��[w.�~~p�(�����ŏ�����3��A�;l�x�{Ux�zg�\ʱ�%�g ���}�O6��B���M_�?Q�������[t0
����PT4a�hڔ���������oF�2rrv�ԛ�㯅^�q���Ǔ�����j��ڼ	��t�HE�ނҫ�J��(@jD�H(]@�H��.U�-�*z��]��7�f��53��䞳���쳟��uW��E<��J%�И����rC%6dA��{�f��1�E�5m���_ד��Y�7�����)��B]g�O�b/��)���yy�&�4bƋ~U�Hs��uE��inl(���L�jt��`��N��ht��n�P����W���a�雥w�~�JV:���m;%�mB"���R ��{=߾�,���r����7����c�V�,kC�rw(*�e���#���v�F֜�
���^	��g�?:bu��;&Ism�U�f�Tf�fZ|�]ay X�3����>���޹���Ns<�H�d�@�m�s��Ϻ>���|�~���i�5%�s�hc�k?T�v���eH�N\�0ְ�[�im������6L�!�$,Z��ɋ�f�V06}��S	��3�,�q',���:��jģ��#���J��?j>3��_B��t��*�h1{�yI	���T�ߏ��2�kJ�"�\O������_�81r�k>=X}�C�)��>J\g�	H-2L��#�`�V�IǟCIqd����!��6����x�X1�8�*���1�dE� ���^���X�J�"��p-�N^��*��%l�_��ʇeo�^�to2<�����uRVs����\�[qO���m�̗��>>2ҿ���P�g>�&�(�_���d�/�Y��0ik	g���)�
<<c���A᎟-��L�����_{��tv�����;�/R%{��^��ף>�U��W�,���"�3d�{�²�?,9�5�Ɏ��
�O��̴�&j�[/�J~���ݏd�-2"�ʌL��#���X\��~�M�W�-r�#࣏Qq���VT"զ���d���h�R9@R���ё��ExDu�u�?�ѠN��9f-''��>�6��Bt z��ӫ�(�
��틮Y�AKE���.���鞲֡��@k�U?V�Zd1�2�$wW�-d�@&�A�\���A���hSI'T��C�x����&�NN������IE4V��J��JD�Pxj�7�8�^[�t���%:��!Q;NO����;��@��X�FQ {�-�w]p8ִ"�f��[mS�jW�l��Y��#��4O�����j��
��g^T�s�Ʋr�u0��7�\�Օs?|��u��������f5�Qt�E���OP^O+TY�k{~4�|
�#㝬��M����p~��HT�e�_��V4����'��g\N���J�|��do���*pNnnL'038GR㆖�s��o������������+/(Rh��z��Z67_21���6��5X�̙�݁�#�y�@D���P1���@���� ���%��a�D	Gwd�EX�)�1�/SMw;�>��Ԋ���=LS��[��P+ d�95� ����Ŭ��z�k�U9'�0KY�hW �Z).Z_��?�h-�D
�BRr��L���q���n:G˦*"���
XSu���%�����nB����o������_�#Da>�A����(h��e��J\,��E��"�ח�>0+��o �#�[�q��B9�Z������ 0䥮W�*�!����;Z��@�:�O�@P�m��y�0� l�#�/�0U�DH�Y�E�_t.#?T{Z�V�L֗��9�1*��;i�0�m�����'�̽�<v�T�ޢ���/4Є�Z���J��Vkf9����FI�T�ԙ]Q�0B��N���{!�6q�vƻ�
��O��C�R8�����Z�	�Hۗ�u|����"BZ頚r��i�v����ɩ�&���`��:c���mK�0 �},��ϖ�8m�|����a�ʳ�'q��$�W�RG2��&���;�|}��� ����r6��J �X�2$�����R<���!V�a��PI���{M�Fu�٫�04��+�\��7� �_Ri����*u����'�Y�,���"�Yp��p~��6vvvi))���S6�2>Lm�w�2���)����2�2R����<S'H�T�d�
lsC5�4��?<�6���`?+�4�(X_�[�l�k�iZq�Jz�V;!z&�+�����m-�2Rl=a����𺵦'S��9R��btuQ�t��9�/u|"lgR'�Z���_�±�+V�8�D�h%\W��乚&�7�mJ$���;#y��O�z^x_ 8��y{���ADa������.��x=���D_��*+T���07�5e:��>N��(�][�˾8��ୗ;D��0�����Y�8����[�˞9�����q��G���b�ǡ��2t6�<т��`����x���v�>R)�k����'���/����#d={��m�Y	~�b#t�h,��.NK�V�+y�YC��.w�NYT�kI��>��E�)�-�gJ�.Q��B:BHG7��n�s�����/^�s�].��;�@�Ҳ��g����Lwr�H}	�1�� 9fC
}@5�}��i^C�^�V���q�#�9�U��a��~�O?�
jw���\��&%��z�	�`�$' u��:�k.^�׹��{��>�_wڦ#*���_��g-Q~Q�2��E������z�m������"�$�S�|�E?�h\���1�z*���.�c]?\]s:k�J�/,P���S3�_�����_�ƪrEB��K��}&sR� )i�Fx-q��N=D����!AEت�il5�Fh�=�[͜/`�k®�xX
���7�0c>-�{��L���[��m;s�S���RHŠYg{�۷��0�������t?�6�n ���X5U����&���n<��u�r�JH3ou�˭wM��r��%<=+7�C�ۮ�Q����rj��T�|��Y)�N���*z���Wz��Ol�}�~6��W�L�2�{����j���(�d�HY0N� ����C�ng"�Ķ��iХ����j*��ZFfl�	�C_��n��A�6�"$5��!�K�1�z��)�;z%�^qj����b�w=��d�W9]��<N��.�,Y�?N�n.������O�"��3�fl�B����.�2*$���T�g̕/�v_J��?�jI,[e��{w-kǿ�p`���t��H�ÖN�p�m�g9܂-F��2��8�b�M��� �ꛗb���չW�'5ԛ�NW�P�̖y��&j����p�7��p85���[r��$8�֔~0NC���H��k쫇a|�yee�1����'F�]+"�x#��zJir��b�u�CS@06��4u�*Y+�	.��'��ƦE�VO����^]�*C�{2#cS<X�Ɔ�j����w&s���Vz��eE�R6X��F5�g�BU�t)۔}��0{�)�&p�,WEP�tɧ���MV$�΍�2u�8�������\��;�1��𫡌f�J� =�ɒ��w3���W;�M�b�*)��H��W~�V�I�5�O�{���;qx��o��P��锃"����	�A���Ch��*�w�Zݭ�^�O\��dx�i5�;ٛo�ہ�q_����Ę�N{�;���h�W.V0�x��"�v*��ʹO�5n�������Y��	/Y,��7���ke��A��ƎW�]�7��/��)f�Z�X	��ɭ��5�"�j����Ki��fY2D5�ۯTm<v��&=ӝA�m����cU���y#�c��8�O{�^w $��l{�@Hh��0�o�k>و~����2gH+[YY=m!��}n��m�7��F[6�D
�Gp�k�/�Z����ܳ��YJr���8U����rwj�b=cyw�i�����qc�˾��?Dpu2��JC��M.��ޭcA惱�ic0_����+�_���b\g6��:_SC.�,���!Q�]''��i�#��n����>i%���L�%-A4�����V^'L��<"\��saw탹��_��>/,^Y`�:��069���Zu�5;[AA��<X�#:��<s�������#c�����W^R���~uV%�O!
�j��K]$�>i�d�U?z^�����Y=�[N�RP�?ٞ���޾�>:�w�Jq�i��	�\b�����������[bbLKU`1`�v��[��z�ּ��\���N3�f�������sۛ����k��V�_(���N�a/i�~mZ��^h�x ���;�7�[��(�4���s�����M�;�g>n���舎�6��(�0���Q,>�/l�HP��!��3ȁ��� 1��}�Oӕ������L�Sp�w��چΩ��HK��r~�_��{tyZ�`�5f���Kw,�(��<C-�ߺ��.:�Ye̲C����D��$Q]^Y1��(�r���Jng��m�"�5�������ۘ�W0�Ǆ��{���_cA��G��xm��g��M{�n��o�6m��ķǊ�o�$�:e~�.6m�k�8f��g�����T��"�U�&�I7,��t��M�n��C�񍤢߷��'���ȘE(���}���jK3L�rk���A��D@���ag�<eD::J�9.]z���%W�֒�O�H�̘�1餛a;�^����5*�W�I'����JR#9�@W86��tz1�B��!��H�9:.�R�`�+���n���L��r8>"G�!��Ǐ2����F�`]�]gQ�4����ɻk�$��o۟X����{�L���./��~���ߙl
�%�������?8`D
l�I։���Yg�8�����RF��U�8�ň���{M�z�6y�vZ��b�X��;e:)I���?=��o���eⳁ��3(�Ţ�$��{��K,W��fw�d���v��@���g�B�s�㙂�tl<QT@;�~7gw�������V����;�� ���lHK���,�TΘ��f, m������,�=f��y����	�I�m����ӂ��Cb��	\?��E����_��ֿ��.{��������Pq/5.�����Z-G?EQ�	1�%�@ �0�):~�w��d�h��#f��Y��4���<fox�D������b�V�"E������&o�E���jT�b\Z������r�]32���E��-�BCp�������&�E<Id}���"Ƴ���6lT��K�z�ļ���;�4�7n\|��[�J�lp���!�AD�x��0Τ/K��歭�­:�8�+]���ɼ���J�Q 2��]��~��
�)���x�`��D�00��8���/p��^��q�ڲNu��[��{-�2��E�j��y��U�J$<+ #�VW=�q�&�Z��Y �6[�{U.Hd����%kve1���.�,z^������%�'���O��7c���H�+��·}��㶞
��ށ˖hj�ӄ#��.o֯tZR|�k�/��)#y�f��'�H@fXs��n�Ш"V��m��*�U�ٌ�~�p',����~:�\?��P���������\+p�gkP���
@�Z	��;��Ջ���@(����d::���)�R/�v��F�6m'\ھGt�q\���3�;��~�0�Dt�ot��t�ԁ���ͯ��q�r�p�M�H�g��d�~���Jf�/#/���a��ebhg;.�N��r��͠���p��޻�$.ζ��NR0\;�hbi�>��T['B���Є"�6!M�SS`��~�(����z(̋�)�Q����D,7G����`���o��JUN�GƦ��`;S�/XOqY|=gr-ѻ�N��!!*qz5�^k��9ĩ[#3(Ʉ[�8�����?b��K�<Q�$Ԟ:B�n��2�Mv�y����c%R�nL�y
�5Z��w�/菑��!/�7*y0���*�:�]������rtŚh$��ܸ�I`N
�K�n֍�t{ᒧ�e2�����K6NrzM;@�-*��ǭb`y�^�G_��[�_�7jj��1B��c���N0�V	���b/A%^9���y	�r�}`�t�w!�C&�|L�y����ߕ*Я:j�O�@0rF������(��R$�dg���x��S�A>���ڄ��y��������:Ij�ih���c���:hJ��Dm��G\���3�=�F��?b�����������Q��d7:XxCj���9N������(�H�-�%���?x�S��^���< eK��q3�%�e�(+��P>=zs�E�7Y������,�P��P�Y�*��2J�~��DaT�=Yb�m�ű��������� �(6Q«�י?�싴yް�[�˒Q��<ojoh���P���o,����!x��E��k�o1s�n���m�&ry��;s�KZ��"P׶���2UK�7,��.�~�&˫�I qs�QOV�����)�F������;���51���[�G�������6��Џ?��i�W�~/��%������~�,�6pus���fY�	:"�jl�7���7ǈͻ��G�������.���ً���<����`ff@�����!�G[!��� �t�lοi�إ��C�8e�6��g+G "�� N��W��d ��i 0 `M���i�E����n�mԄ .g���w�e�� � ��u����3 �\�Nˑ!�/{ĭ3S@3/�T�T�~������`�E0fi�ׁ�~�гF�6ZV ����|h��xuۙ��; x?S�n�O+d�%hX(�U �
=��]�A���b�
���W���+��
`y��%7�؉������"H��\���V_pOCf���JNoK�!��ED�Q��2�j��z��w�h�|��O�ue�և·�=?[�UC�R�r�=�a��+�.'

�Oߧ�A�>�������+&�����D�C�+1�\֩%�������ww�G���G>���_og���������;��D�큸����������޳����U�n?�/PK   $xX~��a� ٮ /   images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.png\\\S�� Áh���P%�lٲ�LX��,��
BX�Q���%�A@�� �0Leʎ�gb!��b�����p�=��y�sB��#=�=�{ /��E���-��|��@�W�]~�a�<����7x��粅"������	��Q�K��&�����N
%�����p��I���%e^S����iP��`ȓ��P�ej�l�{�y�o�!O!rݢY��بߚ愳����}���r�Wk괡XY?�q�?�üh���!͵�/V��xt�e~fc��	�O��D�:���s��;%!�E.�o���˘��P\hV��rɘ �;����TS��{k����EA�n�Z��2���|��k$8V�p�N���$&��������Q�9�HO�	��T�{���M�*��o��f���̑��M�<�!�f(nQ����P/ h�fvh̜�,`�*�Kp��e�Wc=W*&���s#�pSx���]jr������Y�]`7�핮��jʿ#˰?!!�\Y0jn��D� ���Ȳ���h��87Mr�q|h㡴@~�K���g
�	��Xy6\���J��ځ�ӏ�u#H�u!�}��K�����%%%v�ou�V'���'���$�
����vv:o��Dz����p��r��gD�*������Tc����u&�17Jw-16������p%�8Ec��Nl�B�{Eُ��^�LG4� �s3�Y&Gބ0�F�٨����?l�HIƾ�䦚 Y��q
؜$ȁ�,S���fDz|�e,�q��傆��Vn����@>$2�r$t-�Q����a��o!KʐĦ���H9�mb�����m�Ž�u_���is��=ۚ����1�r�|ϐ�B-a9~X
j�MD��+	��#ҍ�֘	��1//�����")�	p[�e�5���(ۯ�N3�� d�)T�����ɂ:�x�f�h/G���%�����	L�e���fx{���}~~~��J�1Ε6/c�&�
?LDD�˓��3�{����g?�eB���Qsn>��>�2�+Ȯ�\\�1%^�+���q��>�n���R6��]�]z�}B�u\����uv�Y��H/$�W3�
&d��Z��v���#����ї����k̉�����ڱGw4ʂ��W/��� Ɖ��OP��m�*�E"7f�TU�����a�@���+���=�o�a5sTL̖=),�Ek�k�:V�[o�_�#� �zbўׯ�o��Z�Wud��x��CU/��Z��,L�s�ŉ�kY�����"NN�9�s?���ma�����i�-g�1����H$_g���d#0[��n�����S�Y� ���>snBj���ݗqt2�0�׏�΁J�����7Z�|�2��_���R�t��� p��Sй9;��q`;6����@��VhS���[�0��o��V�e�_|B���l\�Qq���So��D�����[�m�~��B��D,|x*.F�Ƭ_�8��J$�Asp�y�f
<�]U6��Ka����n�����#	,�~��=w'H�g`��w�z�<s��@���Y�Y��F���#����e^w ^*����&���'�
o��$5�8����j�����	^�,-�%z�h���K`�kʋ��Z��**����J`�W	����5��#��i���h!����6Q�#l\Q�¾��%I�>}����t�=y�y��~pyĒ;�H�Xc�u���޽{ͨv! C'����|SE��u@��;�u6.^��~pG��
� �ژ�m�@[�:�������EEE����G������b?�*���������6��7)%�iv֣j�kP~�Ӑ.�Ă���:�tD�B|{B�B��Ǭ�A���*�m^Y	R���_
�~�VP@���1���(g���l����ˤ�E��m6����@��:9߹���п�YL	�i:��fdZ�c�Z-Eջuee�KY]���mUCEUUF�VT����206.���J޲DvM�d�|�v�3l/��i���9����ϴ��Yy���3�;ǲ���9����vnHa��zC���d�?�{w~��|2����r��,D@���ͫ�P�[�kᅠ�,1z3��@Sd��o�<��Z�x��Ey��(韤�����H@n��̮��0���k���TM����PSc���q�h��m(�Y�
-!��a�؄c�o{�����;Ϫ lv�R�
�eXR9N��6��c�ݽ�j�y묬,�/����bF�a���؉����7��Bl=h����>�n��P�J$�\@���P�y�m����_g.$%'7JTc�e�NLִ����������=�g�'?6�L��U��N��=��g�j4B�- %�O��@%���7U+D���oM�"\�"$�p�� {��+#1���G��P������G�8�f^U� �!߆P��ɲ=�Lb�ض�>6ʎ5��-�m��X�7�E��EvQ�K����(�����- E��ռ�*���к�01>�s��� ')���.Nb��̔�98�p@��b���w�X ~*lD���w��-����B�@�=v,Wc��=�M//Y�o�+����R�U���^_�&�}0sD6�h�I#ql]E"k�뾤�bS�4�]��IU�l[�I��^�7���z�5M�뱂��@��l�wTh���8�4i=8�j|�ߛ�8I��
��$�
�}�{<ڄ�o7�C�+S�$�qU#�3�FFF�����r��ၞ�Wz1��c�N�M�cQ����}�".��O����*m��A_��o
GϚ х�ie	+��dH����Q�kE=$��m�2�0E��趖�`;���8�31J���̧(3�ۅ���w���J/�:��K�\��"��PGe�m��=,����Cj!��W�cVXU��L||*�'d@��������Z�2_9�^uj�B�.+��!1���RݡY����)�&)>�B�פ��HkU��k`"�c�/�oS"���ʦ��6C,��x`����vb^�p�`�Q�Ǔ\lsDY�x�,P/}��r�-i���Y���5dx�w8���t���6�#�q�n:��������f�de��=�����Ĥ6)3=A��\&�x(�EE�f�z�����FWG�l�2�����0�㥒���E�i�^��QV^*S� B��Uqк����P�zK�'T��I|���	Tb�&��S����<��51��W�H$5��(�>nV��*
x�Nh��@�/DDD�$n�'5!����<y`3����l/`���O-P�>��-4�һ�e�U|�\�
�-<idd���v�Çw�����<��[��Fj�f��������L��Ӭ�\�:a���E��)hȵ��Չa���J-���`�[0,�)����
\[��&�,5U�����JT��;6�6	)���/�^�� ��gz�s������]��`w
Q���J�����>abA��V���rkʳg�)��:�����wL�^����6�� TT��B�b���9p٫u��ۭl���2��C�uX���_#	���ڴ������c0�N�����{�����J�H�(�aԏ�Ƥ[����ϧ� T���n.I������;�F)rh���bi�
�Cܝ�޽ks��qF�G��W��9�o/�W�Rm�F������'�m�(&�M�h��z�4�0��z�n�<A���(o���]��4����a�<�$@�V ��om���Ź����+X��H��ޜ��P���~P#ʸe 7�v/��k�4Tj��gߝ���8D>a.�`aiY58ƌoP��UO3���f�ח��/K�j�n*�{�� �@Bv��πn����w-9�E�mL����S��0��/.���WN��_��H�&X����Hnz:�:;CσT�����ׯ_����ۧ��V����K�G�۹��K��>-���f懧o�v5�h>@��'3�a������f�ֽk�mv�G<�S>s�С�xĪ���J�Z��M��k𙅅�)����6 s���1K�^��@�z��ʵ�*�P������"7�rͽ����S���q͹!5`*�/Nu�n8�+��4`�0>֤?<������[+�/�?^\{�9�F㾲�N�R�������d��Ҳq}-kS���sֶ&t�ߟ���N rMJM��Q(:]|��}J[��r+�G�	]�E��]\�JlJ����5��2���o+���T���|�j�R��F�Q����v�\x���%cn&�'l�nP܉��X��М`��C�����Mq�ي�@hz�`�KЪ�,��Y�{�III�2̭mlFD����g�*,�3�=3�X�ؠ��i�y��0I�����P�0�v��qUI��.zn�p�f ��a㬉h59�f�~�P�`(�	��D������,J�`Y��G���T �a���c�7NY�{��S�;�e����3lgL� �s{N�>����$�5NN�Y�%@X��E��A�L�`��``` }����?}��xWt,		��8�
`;��	,���NM��W�^��	�`��v_[��xK���Z�
Y����W���eƒ�@�;���+X�\��XfyTX���C�꼩�o�gwk��oS��I�/����ơo��Y��Ü"1�<�"Q���_�|^�����TSZf{K���kEӌ�'�2j-o����������n�9��ھ��(M=�%#T�c��
V��%�!0ܲ�ܜn�*�ӛ�|�`Y��� ֓�Y�?��-S	�t�&r�K11R�Q֊ ���V )P�L`�����tn�O�֏�#K��bmY���Wy��`�:��#֌mpE銰ʗ��1�!'+�i���>��Y��tT���@�`"k[��%�2����0�nG��L \X�x5���u��4�3 V��`h[�V�L�ri�{K�Q~�E�1\�7�LykMU��+ �Z0��tʷg\Ē�ءj}	DrL�45SY��]�i������B�,B5x�s|�����5�!	����jz���?���m������	�X���2�JF�Vh��>���`靵�_X]��f%��}vu��o $�}���6��r5q /,�Fy��N���<a�
���xS�K��4  \�C5��r��/7|f�}�U���ɞz���Z���Y[�]_�ե ��߿GIlMȌ�p@〩L_�0��r��џ<M��}ZV��5RO8�t��.�@�w&E�_X�Z�T�,,\[����@�W���M@稠`Uy���7����h�b�S?��G��B9����~�e7��@�)���������]s��a��Z�u�z�$�{��$3$�����COh����ۦ���i#p���&J�!�;�\���f?i������E��M�gj��7�OH��d�rйN �`?�Z��x�%)[;�n`����O7=����޵��Ngg��_6���~�rq��'&ZӚ@S�N~|�8&�v�'��c]��K�W��1��4r�	�\<7��Z���߯�>��X���IFݯ�mۿ�l�.k;���!	� }	��3�zr�{��]�"p���2X]3����5�N���K��-��ɩ�[k`�Nͬ2�PXo*���r�y��P��M�A�Sk@��=d���*�D.��'{�Hl,��A�� *��.=�zs0̑�e�oQaO2@���U��o�,� N�wG��Q�'V_{s̰�Ƀ���6�⥒ң��������6�@ث����#|pI�e�(��	8k_�g���C-tտ6<�'�W_�p�ڡ���YAM��&�jSب��}�_J烜��X���l���S�n�%� bSk�P�1ߟ �he��X����<��7? ա�8��J���X����k��<^㲭i"��۱���S�A�M�T#rrr�D ?ы�\g~�(QQ�fV��O%���,6腟g��K`��<���s90���4X?�B=����/,���~�2y�a�[�� /Wל���!UY6y~ڴ���4$�J������u�g���W�}�8Q;^rݹ���%ǟoO�z���U�}�:[$�p���y쓣<��bmi ��������?�m�-O+�T�X�������u�2�xs`p?@�C �c��B�R�m`��0<ˏs,O�V�x�$�C����c�'V��[S-��K3�k?>�Q#ǧh��8~qnC6�������\K2�L�h��X��ꇶ�˓�C��Z�ִ-��@�Z�E�Y�v�5��1�ָ+��-��ָ����%��E�s��&��s/��� �mqwb�X�����|a�~ds�g{�B�DA{Q�Sqc������D�]���Z��,�)��y�X�O�-��<�շ$׏�i5��ʡ`,\�87�Z���n��`j�\�N��.��o���E�����{�ID�$6��!�?/"6{���a0Y�*�v��_:��ء���~�.��۠f��a�c���B5�:��ڶd� m��V�d������/��R�й	�����/P[uC걣���\Ǣ�H6�e�ϫ�J�PuףF�(#Fk�l��� ca��/x�����&�=��r���3�!uQ���{����J�>Q�ġz�h���I_+�1�L���C
�A�h��C��\m�&�O�j��P'�uE��)��a���������˾�ޡ��r��SbƢQ2�1S��ݐs�;n��D�m�Nw2G�Y�!ayO�O����dY,C~U��!z[��K�����p�<ۋ�|ܯ+��0�gϨ��m�az�	���5�{�RMY� �$�lz`tr0�f�� �G�v�V����:�_���Ƚ]�wC
������r��T^n�Q'���n-�xM�$�����q>!^�h9Q��c�@nא
�Ճl�n�_D�/�����g�k�a�2b��b\�4� �?�e�N맃E�D+����0�j3F��
vz�A*_���p�\�y�;o2nt��.x�9�qAa���}�1��J��
u����$��&ɾ?q�h���}Mؔ���2�����۬$j�_�[��A(�;,��+��I�7��A�Y��m���++�O��,�$�d�����ȡUFH��(�S��:U���w������!0��FͻL�5�=�g��vx^_�Jv���>e�b��Lg�V<=_�8��h��>y�0���61���j�O_��������@�X�p�:I�2�qm�/�}��RT`z7���[�a��V�bSL6��ˆҷ8��7�WUH�]t�PI��)c�1ùw}`��[��9j�:@����1h����[3d�����{"4c2/n�j��;�aw�L,a�p�`����y��C��c�kT$y��3�����8�:jR��e�	��g����`t9
׵=T��
H�w⨟(3֧��������Ĵ�1�Q&�m������߁sHw�7��1�	mK�m^����Z��rA�y��+H�b��j,NO�n�"Į�HJ����s�d��!}/��6�Š_@u��4 ��w��(μ�4��Ѻ�#*���t,0vRd�8ǗC7!�v��>�S7�ǤʑA\I�3?Y���H��U�y�&�v� ʴ�i[bp����;�E:��:Z#&��a�ua�W1ߒ��HUY����ˁb��D8�_��W��e�����eGL8_%���ȉ1�$oWu;B
�?�a��tT���Xm���ޮ��:K�pg�����$̺�w���!��vz<�:KΎE+��j����qj�}J;J8Y�r����B��t��:BS߼��?_�Jt�vMtGF,�*,C�p�G$]�	)���ȵH�͟�O����!KOz�ۤ�Wwzn_)W?(�OG��>-I{�N�)U:�a���;i�l�jw^�/�VCA�]��%�W�g ��/ӟB3��7`DsL�$9�U���er���4`փ1&��Q旗�<$�1�3��`.\e(��:��*���C���3��ѧ���"����N���=؍��%κ��
+R��8��čA�.���2�p8�Zo��tO�v�h. =X��	;�^X������`��G��v�����e�3&F@1���`�������A��;D��0m$�0������/�z�}��&���60յ�� o�v�O�*%�A��ݳ�bz��K�v^a#e2h�8j�O��`+��9�v����O�&� ���T� oA��&G 7;����ϒ�H���ə�Ab_@̏�h����J���/�R 4lg>����Xкщ���̋0KV���.�b�����OF/z��B�]��#v^��1�3�8N�N���i^������xЭ2��dE�+�v����@ƨ�(����H����L>����g9W�1�=��i�Ϯ��o�-M2��L�+uw�6bGj�� ���g!�۽���N�����#��h���!Q�!��w:'�ea��Gb�YP<���W���<���j'���@��c\��uŚ_ND(_�y�[&�O�b֯��p�9���-���´�1�7`�]'x"Rv"P�N(,�d�%��,9 ����(G �XM3�\�����H�;X���Z�ť����>l�W���y���?+͇^��)χ��?y�9}e�yZ�X��$��c�i� �S��Mi�}6~�A�)�����qh����!I)���	�1���9,L�<lL�@"��8�~Q� )vdd�*��2k�Aɀ�p��H��SG�����!���p�M�1��Q,SHCl�P��x��^�tG��_�6��5Ka�b��`� d���/���y�L
,P���0X��N�K�bg�u�B��Ǝ��D�������G�Mc+݅����8#�o�&�25D������jV~b�u�3?y��������$kY��y(��G�01����u���hA�0~l�����ql�ߤMݑ9��2$"�s�h�]N?���D���Z�#��������D��k�:�8j�yۏm��([y�d������]��z�����ioxԐ��D�6/aj�Dk�� �_f�/SFM���l��s	�ߐ�C	�C��v����V���2��5��S�|�����XX5tNGŮ��SE �O[mC5=����	1�n�G&�ô�{���WN� ����'$���o)?�QXH82y���g_k��+��vG�������߂{�=-/���fk<>�d�Obnn!_}����o��r���-�rl�����d��p[O
���kz�����P�W�/\�-�=~��4r�=��_������?�|y�TJb.��H�p�)k�z���i� �=Pأ�l�f�����(ͷ��)p�?j���{��۰<�j����ϡ��צ�g0������\��
� �|��a�b0��\�;,ƕ��8�s��'7��szr�ߞ�M6��>*�6� B��<��9i�N�}��u�	�%�ﮦ���%Cs���$�Qҧ��jm(&Ց�L٩fl=l���8��;ҾlMi����W�M���E+�zp���� �?2��摕2�����[-�Ӯ�_����B�{���W]}����E�H��e{���k��>5]�i�W*>��H�P��ݭ�G)TD>c��R*�����#�ɐ�~A�Wr�͸�x�_t���T4�/�׈v�����Ԁ)7�Lo唏8-"?Xͩ����o���k�w�'�y$2�����,�����Z�b�ٌ%ņ:��s�N�g�)Ƒ����(1�M��ɘ���Z�q�q�EA��{�a�}Y��S>�+}ͷTB�(��T��"�&�Ά��}6��>�}�;�JH}�[{�(�ϣ���%���[��!v�j��(��Y��__t?��;Xȱ"wp�+���3����kֶ0Bm�0����1���q2���@�����I��g3�"�^�NTŝ��������0ب���U�0D���7���aK�F�罹����g�+5j^��q=|;G�= -{�BY"͜B�ή%�,����^��o�l��I��HF2��-1˭�]����=�o����}D}7�����a�߹D0�WЍ�0ą��%F�9�2�$�ך�:h|%�y2������rYHJ����ڌ�)�鄲�|)c�쳻6�8'p!q[V׃=E�;L��K�Hi����Y�G���:��[^G#Z!)���Z�@8lE �^��r��ݼ�C��4}U@#H��*���Щ���W �"H���v+`�T"���/�3���8H D���p���ri�-h����A�� ��4<�X���k�0���u��A�]�<>J�����3ag'2��� �����V>����߯��m�&)�Q�H��r�L��� �g��;=�РS,S^��8Sg�u�G&B
 ��o�d[^�=�+�[z =��{���e�ο�Wj��fa%�>���ɴ��ڜ��i�*zC���Þ�x���Y�o�75&����];�:�
�ŵ.MS<�ͻ��5Lh��M�vi>N��ﲽ J��O�+[�¢θ�*�7�z���yv�%��a����Ӝ�P��Ϻؔ5����~��MDɽ!� ��0����~li���u	Z�AmȀ�sV_���q^���O����N��J3���#��m�؊2�!���FA�n>��N���df�)|z�<�>>��$��"rO���M%���&s���32�1�=Ј�����Os׿���v�ushD4�x<����H����:������-m�S-/M�/I�
�szq���f�@�M��X���bczg^C�:��/�����ʮ�]�f��0����U�	vmCѼU���D�U�� �v�2~��O�ē��ǡ��.���(銎�����hкL�_�U�်�G����^Q�O��(�pT�����]rf�	��Y�)CG���\�MON�&��U�Q=��ݯ_�C���>�.�p5)=�98X}N�󮺺z��R�vF�nC���U�lՀk��I��p�u7�u� ���FS_V�!Ô��so>==ݰ�Z��9��E����b�F��<�%���Q�W�W���f֝NlRް�E��.��ux����o�ᝨ�E-���o8-� ���t"~?���jDJ�D�qU����'������+���#0�3ٜ��zz޼'ѯ�|_�H��uN�������T���kB�(�PiӕCU��3)_ߺ��^��93���X����ٳ˞�����4�k�}����!ct�����1]�/6�a)��R��~�ʸw`��x���'/���.�����xe�n�miӓ�'999Y�$����7�/!6������N��8� !��̤�%�u�����y^�6��YNWE� v������jЎS8���dwGxCPl�Ӿ�˖����̳�u��8�3�[y��Ŵ�͛|��G�$��W�X��,�����ҥc�G�ʌѱ$F��F��,���ʙx�!36�D��gm>�t>���~��bFb)Ԇ}�kY����H +K�ԇ?���@%�@������D����-h��E�>��psE���"1ؒ��v+�����	�,�_`��/М!��h[5W�=x~��	�Oќ$��l�9�:"�Exl\���^���kV���o��l��:���y��8�G搯���3�9� U>W�٘�'#�>/>I��2��{>T��I��!�aBV�c�}��|�PݯIG�Q�Hk��Ʃx���=����h��������Q޷N�m�i�}���~��Ec5��ƍ��"R�?�˶����uO5�@li�4��oyL�Dʦ�vJK����9nF�[��{e)ڕ��������Y��3q]ۺN���͹�WD��
����X��̺W����լ�
�{�����+����3�cqM�b�q�[�o�}B��Ç�}N�&b�����7�Ż��8�+J@+��g�� l�s<�}y�=�Ϸf*�;:�<1�~?�*�)��$��,��(l��P=6�<n�kk��<	.
G}+�=�Μa}L�]���ށd1�!��n�>̪�s���>o��2h$MD���Dj�׾)	�k��o��?)�$Bd-�?ݢWg@b.�t�|�!:�t�	t*��L��s���Q��$f�79��&B��$&�4�6*�uZp*^`�M��)��aa�	�Esqǟ���β�J�vp�T!o��#�'h!����ğ�$��]���М��"?��-��k9`���q�����BeG�K+_(��8�����cxY>��1�O���Op ٘�W�b�PS���Vz����U�oj��uU�.�c4���sw{.ތN	��m$]����r�~�z�L����|�uM�e��u*��<O������L��11�H�3A�mUcz���HʎH����co��m�8�3��.�>{i��/�p���7��Կ�DL]�EtP]]$i���Pl`ĂA�u�����ԗOE\OJ\r�nN�byZB����\����Z��CS��sKh��9l���3�^jn�?�\���,#�Dz�#��Z`�'nPBI�S�K�'dRo�l��j`I-X�j�7�3>�[_ooR�n"ayI~.�%�����RNhe�3$@`�O�k�Z4/r gyt%Dr�Wf���׻(�,�VMryqE�&�}�{(����	����' B��^\��{8YH�[�$_Hf�{?��c�R�kL������0�F'��s������NIF���\{�����<�˖}�s��U��)W�<-��#��&@�$G(��܍��DP�B[��<��@J]{��T�B����ڢ�#83�镴U�tٷ��"ü�h�ZyCv=fӈ�5M���hő�ˋ���mӋ���/:uޓ+"2��PP6[ͅc[8�e�����>�~�������δ>>ӢEP2��|�7�w�k�
�}ө�y�p,���S�<����R��ܛj������w��_�T�B6�tH鷿[�XEx_\yų%UN��]� guv�_���4C��φ��o��Lm��U�)�@�D��d+x%������b��"@�lv�����IR�;d��!���^�����In�B��4i��S�6w3���x#����U�OTG0�Wწ��;88H�U.(U��k��搸�Ǟ�����l���k��sY؄@�1�*�J�R��^�"�/���2��:����5��p؇�M;(kH�������d^���/b0ݙs?Z<�Ry- ���������Ч�����Qw��Q���ޙV����I5$������+�%g�S�b���n��~�qe�(淞�*�ȗ,��!;R�ҿێȕHl206�XX 8Q���1��c�T5nӡ���ȦR�*��SӔj����:0����hI��2$K��$�N���>t��)��Sq����۷��={��u�q�)��~��%������=1��)�I��xS� G�-�?��pN��Ԗ�����4���,
��-�r�1=u�g���lC�}��E�u�ԃ�G7��i27��cҎ�{��Y���Q��&̚kW��ێ)�4]��E�{`Z=ǖ�{�7�NI��X2�·��D��t<H����%v�~�^�����S������ �X�v!4�T����c�#���4�-c�j��3�ʗ�bO֯<.��dT�DW�h�ة2��Ə
g�����=|��|�����l��|Y111A���n{�B�ȱc����Wz1b��j&��"H������,մ��`���Q���6B
�t���Kk;K#'9x}�Ћ�/�M�t��/��I�N	��xC&�Aȼ䪲��zZ��Vr��7����u�h��n����(������G���z=ο8geulnn��W]�>���422b`d���+27�,��I�5�-��8��[��K�8z�͹�-Ȱ��+�w�mS��l>ϣ*G]���-LNM��l�����L��Ż�����}�J�Q�n���:�d8j(�C�c��P����-��-=�% ���<YAJ�t7�݇V|��V{���߄)=�5 ���[8���|����]��G��Y���@���'�kJ��텅���r�t�(��[�| �
��:}j=��e��$�;��g&ք�[��?*
Cph�UK�UK�j.㯜��b֎r�7���}!Dp��
�R6O7�M�k �b�Z��9���1�{1��	���@*gخ
Π���3�}�iڔ����h/ |`S�,�o��L(][v��;8�J.�e�ށ��1_;�1��f�F��6Θ#����&�氯^�����t\#�qQ�|�8���Z�.������R.?�vY,V�7M�d|��S�5�C�M2^cb0���Gu_����d�Ӈ��F"�bccn�K|���_��f�U�V%E4�M�� �"��$������6VI1���|w�Zk��`Ւ ��Ix�F�#�}���m竾wa\����ڃ޵�y�!���dn �-�ڴ����@��=�p��al�n�������O��R(NO����[���=
m,SM�>���ܯ���.Z׍��:<q)o$�8�PTW_m?2��j'�y:;;�}�c���7_(o�z}2gI��s��Z�ZK�|�"�|(�^:�to�+�LK�?��tlJ�)0*<�l�eڻ�y�Xd�35Y�J~Rc� ��~Z�U��(o4lA5���\��G��)��$cX
!�����W���z���͑�G�U�%e����[+�ؔ%�.�}��X������VO�-�N6Q$�=�0�Qݩ��乸��;������� ���@TҨPu]к%vU�e s�I�p?�7Y&�*%��fL8 �e�^�6�����o�2��=I�Mxw<�7&��{��8Bҕ���^4�����<���/F3�8[;i��t�8k��P���P�K�����-����ص�<׿V�;{��; ��y^�՛�Gss	�U��MdM0�{����u�|��<�;v>�=�Wy��,����oyY[�n1uݼ�v�Y��	`��uCa�:R e�t��X�M���\Ȗw1�&6���[�����|fT)�JV��z�6΅��̱���%_��\���s�Yw�$����sz�������;R�UKi{� ���4Dt'����� ;(���*# ������FMf��o�z�0=���wz���}x��`���w[�|��xOrƥ������0��5s��D�1���rϦ����8��zR�⍺=���~f���[��� 5Wx���Ytmk)A���wK>���V3W�O|f$L�XD[9�������{��l^uҋT�Ƚ�CH���k�B؈Ɂ��.A��L�>bhH�Xl��]��ݟyް��D��O�(�^�Y��~�]���c���֯��%��e ����{翼Ɉ�/FQm5����'�$�``���1�ɽ��|�,�t�@������9�\g���h[� ��d���3k�yJ��D�"N���u��$+ל�T���LF��I3	�Ћ2\\�{i-ۣ��9��7�	��-ة�����t�q�ri
]�"A�ȹ&�c���`���`胭#=��O���T�=���0����M��#:)dǰ[���#�V�T>a~�Ź�#��m�)�	�{-O�ݬl�!�0��R,�N���ʙ+��`��w;t��.[���ϯ�h*(���((�}rr2tI�*�@̯�����JG};�����>�M#\�s�p��m��7 �-}?��vgؽFtm���D�쒋�3��ߢ*�Gt�����g�}��_��lՃ�=��Z�.��}�ֆ+����ߏ��mgv����7F�\H�@���n�{-05�N���I<��D�q8�7چj��r���1�9tD�s@��@�����q��SXӧ�i�H?+�~�����T��������<�J�"sM�;Q�|��YY�#d��.`������9�����`m�*g��ܑ9�UZw}�>���][0ӽ�yW�J��ִZ�u�<jӘ�o�.I�n�y*#l�<�&�V����9�L������1���.������7j N[�S��@��myfw��J�G�@���EF#�3����w�ҋ\{��5�J)|��;��'����K5�W��4��: j������F��	�I�?�jP��I�3yb��i����=`����/�>� ����=N��`��=ϓ-�4�����g먬��43�8ywA�뵳o��C��g@��� ��5ꔼK����8��qV�����o߾������>D5t�����R�e�Z����3���kI�sW��Ԛ�m\S`�Oف�(���1qq�CFY;t?ۖh�-����	B6q�ޑ��˨�vZ����S�G�� 3�TVF,�r:�1Q�������]����O��X�,�,�o��aٮ�ȇ����V�5]^�1q���!2=��S�<�z��m��jz����>��~� �G�qh>�u���}�j8�q	��2Qb��x�����^�c	�f\�&���lPI~!)O��m�~lW�KL��� d����g���\�����Mw��Qr,z�j���5�X�QAAvʿi.u�H���+)��� (J��CL��h�摊��59���S�@��000������]�wo��^�=���<�0�4hF�U�IѶ��n�6-�?��8��W�_7���D"l>��z_���XZZ�q�gb�y������=�v�c�Ho�J)%��9��$�?~�/�XDƮ�X9}�	�]@����.�����xY����r-[�eB�d�ۍ_��+F��]N:q"���o������ֲz�a��?�����Mֲ���U%�M���t�*!H<���ag�  A���ޒSS�ǚ�Xᣇ�lu!�.��N�*$5OQ�J�V8>�es����v�j��< �E8/9LA��-��>V!��M�~��߻v�ĵ�$��rv�r��$ Odyy9hy#̗�/NF�������Ϯ|��t�3 J<"�f竾�	�a��+1 {��oY?�$��$�Ν/u|�����U����}��0�����׾���u);U�%�)*::L�~�ڞ�Jw�zj?��Xc��p����S��9oo9�ȰT�|��Zeo�����%�d�qL�B�w�b��sm=�:�a��JX�;ݞXz�3{#�Zs::: *|F?�>����8��7h�ug��Yڥ�#�p�ͫz��hh�=����-rh�:����wU.~qcmMp��8�E�D]�А���m�?Y��Xp��M@C�p/�cmPd��-;-�bd�Y��rH���+��[��R8d�g��YB��$[8[�&�~�2�xN��x��N�<�ԇ�C��{}y�, t��ݞ��"�HK���嘪�h�{��?R��>>O��U���LLL@n  ZsL����I�N���J`�VI��u|����ś�}��|��~��3y����4}w<������HV��Q�){o�P�̮d�ۑU$:V�)#d��1�DI����>N�ؿ�����q�sw�u����9����K��۷o+�c����jxԝ���^��j���mO7�*��&Db}	A� ��'���l����Ȯ��Ȇ�_�i��9��	��.�7��H��h���R��ǌY��b@��zM4��Rʬ�S�&:�:���)��qb��O��Ƀ��>�d�r���3_4~��
���J�j
�
�7b=$��ĥ^�: ��,R-�S�9�+]6�s�0}o�h���r���g��X�+�5D@"&���)���ʎ$�����4��G��z�w��"d_�~M�r�xH"Le*���Y��[���-�Ժ�x��Kz��ri���������{.�Ba�7R�⩣u<u6���7���ɸ��No��6��0�0�<�X��MZ>�a�(
��Ȋ��2������N����P̼;�c��a�o��/��HXy)y|s���=�d��	�VU�K��X��-xWX3i C	m��i$	PW��dI�CF�F@����Y	�}�F%���:Н�*���&�m����|-�~�a�g�B �=�2}}`���M�^����0Raa�=Ț�pl��WͭF�8�ח��lh���h�Z��R�؉dg��S��]}}u�)r���e�s������6�!�M�f��ք�T��X���0.@z�`����1���0v�ҵ�2���T����j˶����SW���"N��P���S��A�k��z������;��謽��e�)��
v��$��-^",nG��TK�Dw��8ϝ��M?L<���A@*i��=1f%��%r�]W��@Zk�G
�:���F>�=K�!�J,t�.SN���:��U-��#��/:�F�n_�񵛮'N�ɱ���V1�P�Y�iW�۩��_Қ86A�\.'�=xU! ��N����g\��I���T��:�:�ם��_�#� P�e%�`���A�?Ra�3�P�- h�4d��Fg�KS�y��^j�#19��=�R���8�d� ���{^�m_��3�$�c�|�zu��7���C�*wBBT�aůݰ�21XY=NV�\�L��%Aqpi�gV���'�n�"vK�����嵵��ű�z޿��4�W~�jjf�d�l��m��7�E|��0� m<<*l�h#�,�kkS������E��ݱ�P�nn������7�sQ�(��Z�ݥ�\�TV����Ѕ���((*���<j�a߲l�p3|
4�ň������=&��yyy_fY�9>����<<��9kSO�|i�%�����w�G�K_;��f�L)b���Z-������c"bq��e�Qܐ]�-�!����ֹ�L�α:�%k
�O�kg��K��XX@�O�\�=8hȚ7|�R�htՌ�H�)����w=}(�G�>�V�;A�����w����bꕦ�����K[A���s��!?ޤ��)Y-H�l/w)=F��B��k�����;=�cn����N@���
�̋_jkISk%�Y�ѹ���7Qi���:1���Η��T<?{E���U����٢��v����Dh� ��oݙ�+�T<�������BXbB<@#�LG�$
�|�yt��8��j?1�e|Z@��~����CK�Zh���t_jl���т���[5u=0 �����h�usVK˭1s�5g��x���c�����\�2�ՒH�������w������^��~���X�������TknPbecc�l#v�a��$��7���1�� A%����C<^���	X����\dGG��u=��M{��^�&_�yQ��y�e�`ޥ���qmZ_Ta��zp��2��{s���A=��Y����%���Ö�/NB󌽩�i�K�&�P�Y�3ƹ���4�C1�W�!2�ٚ�T�K-;��x�qq��x���Qw�4������hσT/��@�G�8rz#K���qo���o��A��8���{�v�LF�"�'����]Avtv�J���y����.��H���x���(٢�M%�[�F��E���$+5�΅��kK-h&��V|�����+�R_m�i�)Nω���(̉����>>�<0 ��ׁ��P�(_���rTn�9�J2�IDs1��'6A�N���iLqޫׯ����B��z֝���.��7@��݋���x-y<<�D�kg�Z�}UUb��	�k�����	8�V\H��OLgI5hb�L�Qw`�j���P0�6��c$��7[���Ν?��l�����-%6�8�I�a��	,'[��h���\����/r�ξY����^�SZ_���+�+�D�ٲ�$�K������3��:D���k���?���g{.M���z0&���rO_��$�A+�������)���h�1��0ڲ�G8�n�@����!CP�P( #��R�=��b���y\S9^�~�b�Y��߁&T'�|�G�,z�I�f��Y(��v-��������u��g�4�C���Z��r"��g� �W�V�N���Ъ:��gF�-�~�8��;����z���Jի�ݻv�͠�;���k��H�1��~�{
�p����h���[�-��tQ�w���R��?���vv��|�6Q,�ÿ�����D�7�:w�}��͸흢p�K 
��G�ݎc���4W�t�=���w�Q�P����
���X����ͯ��s8X��B��>�F�����jdC�eb�\]4�ąN��/��Y��`*�s���m�EqR�R��2��f�(4�U\���	P�����x��GQ�
E�m�]D�=��ڀؽ���'i�+��tޙ���ӌ�;��TKK}�����\��gJ��\ZhGy��mv��S�jyd Sd��C�~��!%������.V)��HJ��F�����<.H��z������7��s�^�*�G 9/D���lv<�.�龹�~w���=z���6���%=B����0ۅ��Ҏ��{@��j��慆Z�Ǯ����j�v
Vy׹�>'��5x�EZ�	k�����ޘ�{�T��9���K �G�L�՟RY�
�D4z*4X��xj�5(����7Co��Ih�JN�o��*�����_� ~�R=�e<,�,݃'v`�LB��9����,���-��M���qj ^�~�/������S����?y;J������=&�me�
+������s��k�4�j�f���=������T��t����??���.Pϼ��ԏsZ�b��=��T�՛pZ����*�>��j��܂H�FMo�/��I,j�B�D���"̓BִY���yd�ʛ!ĩ�9���C������cT����⧶8#&�r�P������ڰS�-Y\s�O5q����Ai��$���jn�0�bTl�����ϩ��v��+�nn��3z��/���r-�6ȸ���}�x����꡻�����nMMM�-k���U�<@D��|�r�2w�!lܜS-f;E'����y@���:�R���q��ϯzt�B	L�i&&��8Y��^�]�T'p��^�z��$t��J�=X[�s; ���H�����F'5��B��Ȳ���S�Uq��P�\N�Q٥�TǗ�[������>y�����~��,�������2�wr��/Ma�9_�[���|P�X8-B:lF��_[�ia)'�IVZ��v�nms���� �7��/���2�y@�VTTdV�����s��bU�M��]��c!nݔ �E��5I�^z�R�K�.b��TC"��R+ɺL_]�h�z�+m�w���3���������9 ��9�o�d��+��� �쐏�����D-����G�N�k�V�P��~� K�p��`��l^0ٞ���%i��l�Q���Q�Yyi���mMf��{yAA���w�R�4i��bg�����n��)��q�����-е}'�I�aJ���昹k]��\4B��-�x��ew��?o�w"B쮉	'H�'@m�y�&m�l����~\!�V�������=Y(;w7&��D`Y�T4֎�Dc����!}[Wr���,�>O����ɣs�S���(���ۦȦ>#��:Ew�~�y��g��jڼl"27r\�󗏿*�6.��p?�"��(�,�[�6�d=���P������h4pN��!�y�����-��,�L��`�6�_�֋f��r
��Y�*q��/���(wW4�����&�B�Ȳ0k��шL�ٿfK7�*oߦ���u���B������@�L�_�޽~:�z^l����P��59� ]F,<�C0Rzi��`,&���x"r(���L�A	�	T�5 A��f�#�M�+ܬX�v��x��y)�����X��y�yX6MJ�ib��6L�<���d��ރ�0	Z���b!;���6���ϻ5F^͟�A�GEG��U�n�	r����oR6�ƪ��LD�`>(���b��w���II�m�����鯘Ab@���s]x`�rb�^ʂ�|V~u�� L��z���V����x�Y�����V|\��NP�+sm��]00��J�E�R,AP�(�]�=4@b��&t֒Pj���8^�ؐ"K6n5��_%;��+�LA,������Ä�8A�6iF���R�K����5P�1@��3�o��݌ƙ�B)�ϐ��>Qo@�d�����{CY�+G=�[�GLAAa��حE��Rc��T}
]�VQ6 ���ߚ;�s-���y5;��{�/��E���Q��h�� $�p�f3�jk�����E����k� 9`p��:��$l@4d�is�2���X&>9w����徔1A���ǯ�#�8?�a`^K�2.�i���@ �6�p5�j�bNOM�|�9�7�P��Y��g��8�ݍꍐN/ᘻ�W�_RR��<AE�N8�l�1fn�oj�o)�c#��'���?g<}���dߠ%B�n�[���W��	�Ф�6i�,/�*w����U��/��6CEF�q�3j]\�Ҍ��ܪՕSf��`�нN�� �F�ޫl666�UC2Z��o�˛�<���ߺRµ��� tg��5��<'�I��Qq�#�`P*m����M[�X �� r�V� )�O������l�KuMM����+3=!@B�Q�S.�q�|��'R"(g�Q��i*��;��;l�K8��������g?EtТ|s-:a���K�*��xU��V�0�0���gǬ"`�и����a���ճ�E������)�,S��Iڭնxg*���?4���� �f���Sw��6�~V#Q����VM��,�vq�|t8����<%`a�X��G(�鬓��2�Ɋx��v}ح4�yt�XvO6S%�ӒJJ���[v�X����S1pC�@�K�9����୏VD#
���߾�������C�7Xl:x����9����1��/��28�u�Ctnۂ��P'[`k6�{S�hw!�h����l��YE�C��HލB�˅�3�TH�g^��cC���7���~�8�n��îJ�8�i�ޝ�$�Ey�R��,�@��y����&�����
:쪒�����qR"�^y�M&YN8����4�q͏C��]n![94�d���q5>����V����^�<B��2 ~���*��zWW�J��ZN�����p�� �����KKK�;��Vl׹a���s�YYYP�@&^�o��Ѻ�]����ޫ��=����4QWW!y�Z9��A��uS �#�R 1��o�����9����CIR�{`��f�4�l�6��R'��l�^v�Q�^E8�k���X�1Ԧ��=<,hx�ʽc���A�����P�jk�1��ڃ�A�<������{�1��*,���gs�������ttt�z�ѥ΢�9�������ſQf�[�n�黻>*@����@�����=9>�.�~��W���i7xh�흝L�*�4 �/6�Һ�0���ϗ/2�%fmEF�:��z�\��ϼ��}/n꧳�������T6�����;N 1����??h�6�.�2O-�Qy�ʃC�*F>O�|����º��K-�g�R��	9Gv|(R�2�!F�#�:��2{ՓrS��aS���I(p dr������Z�󎊊����d�kn�����72y�t!�$���1w�B���w�IF�l4�j/zӹ�����)u+h	��z�X����� �`m��/�+���g�.�R%�]�H�������ۺ���ve�i��jӏ���loKὸ���"z�L�"���A������|�H��.��1�}��Y �yݙ,2݁���4̂tvK���� A"4���%y%��v�}|4ʗb&���Qh�o7�����~ỤJ
K��A"7��#D�_ju��h*�>kʤ��[� ���ci����ԤRM/���ա��Lȕ������s 9�a� ��6���f�Loۼ�*?�Dg	�c*�I���I�_3�6�Ղ�������s��m��h6=w���u ���܇V�a���X͝x>���B����@���ܢ�����B�5�2􈑜�:�y�?�43y�/�\��<����!	d��ϫ�Nc?PXĊR���)� �O������T�׳��ӌ���+���\RbƄk�"�"(˟��K��E����eQ��I�
i�?tq�C)B�;���uo����d�O�2���LSts��ؙ*Q�E��W�?��Tf;�W: ��q��Xl}=+={$˃*;Fȝ�*S"��x��.������XkH�픗�w&�J ��x���g���f)��a$�wG��>��A��^�}�|��"#��z>�LW%���$.H���S�cFӤ����]�1�on�p�9*ZJ��6�/7:��}��HO��Q�^o����R�l�[���v)��g��6d�0vO��F�[}y�;�F��C��A�s"�l����K�v�f���{v���h���K���v�C����\�}��F�bI���f%�:�{{�
�L%Ʊ>�{�C�}|R޽{�.�E�ͬ�=�Ī��Ē��e���u-��1��nX�Q��]�h�}�؛Y��|[v!����Q�ˊ���g��:�#jN.Z����ᣒi������^�����9(ం���\��4:'�0���,�~�{��@�m'GV����׹s���?d*���q)>�2
!	�e���ܳ���A��;��Ж[���!K���᥈B=���ez~�z2~.%�y���X�������	=	~g���k'�r(y��VLH����ݠg�����d�O <�Y~J�n��W(��h���v��=�ⶎ�+�p"C`+�G�vy�k

�dn>>�Ý?~�}��5M�[�|��ș���Xrh��$�-��6H�0�4��s||��]Ĝ�_6�|?�D��5G�DV�%��&}�S�D����ZtDY�*�ߤ�x��g�T��SXk�DL�6���9p���v6�������4�$��,�-�]���E,C�(��c�J��u9Taߓ�'H*o[$��P�f�`f�{�@�B�T��NT�j��:oN7Bk0�N�	=����S�ר��[�� �X.�.�:��r�f)K����G���p����ǖ�s���|�k-�ئ���P�_�ʀ	�
?�T�}��%���Gm#��^W4�j�e� u��=��5h��h.5].�条�df��������!@���RC�$�Chjv�
�o�>��P�n��s+��3D������²��Q��!y�2��sՙ�H�TYp��LΌ�g+e���;�+#�i䨕8=I~pBz�1���Y�}��tû���G��$��z���I{zv�:��&zE��h��$���-Ռ���x5��	����
���QQЉ&ҝ�x���W=0���nԝ�ݪ����,��Ʋ<��i�#��B�����[|^ԃ�����<ЈGi:P� ��q���{�$oܨ"��l��9������(^�nrO3�hyKRA��tc��W�w*�R"��@B�EY6�Ю�N��,n��H������A�/���(�r	if�r�P�X����Zw��6�p`�j�*#	a�S�3��N�ц��X/	��?d�CʒC�no�/G-/�"��"���Z�z�$q��+��~=yv+Q�&�=�9 -��s�C����wC��0��c?�Y1��Ձh�����i�c>^Պ\#�Ta3����"3��v|oCd,+�@D�����Tn^����n����Cw�CS���Uk?Gߴ������EN�@Z�ﹲ�(�z��:u:�� �NA�js�q�F�@ΐ����Y�E����8��0����y�UiJ&III}¢���իW�!䝯�}���m�#?�$�oA��	�F��z�̴���z��(����������&���N�s����M�5j^Ck�>��]�M��;���E�~}~��m�Yh?�#�7�%�;qU����g�է!h<d���N7��u��p��,�*mCł���	E�]���'j��{7胸0p�j��8�iEI��w�E�K��Y�7v	f%)��֟a�7o� �g��"�|��Y��7^�<./_h�%����L#p�_�Y�g0�lfG��l׌+�G�{�	"��u����q�-Є6�sr|�ZX�Ub[8*{,�~Be�� 
*֞�+x�N<�xL��Jx�@�����?ڭ�qZp{�D�籋�C���/\�����NY�掣�K��x���zү�X��Ú�u���%)y��[>?j,Y+|NԮ1c�.;��������j���y �9&|~���:wkѯ_�����z�0;�Uyu��4C����٥h&�9`��xAe4�m��/?�Z�C�����tm�]�J��i�mt��{�3� �o��h9׶�Z�9��H֪��l��s��#��"Q��B3w��2Y�xH����0J�K1�����׼�ѫ�F� e��1e�����W�����.RO���G���؞SRQ�k#M ���|�s|�s��p���jzSJ���0��T�����2��ow��H���?�(�1�.p>����KX�J�!�r��D��ۑ�r�?-�l�0K1�o�*t�[��|����&_����Fq�/.��k��g�U��Z�M�������H�r������A�m�=��� �x��$+�]�
�v���XQ$�
�xLSN2Of�b�|)g�����{���ljt�������d�YI�#[%`]�:��S�F��~��p��y=9��#�n��Wh~2��
$ag����hĭv&@^�"��g����b�&bd�͖q;2����0Y���%=H�v����|�G
�a��|W+���r�>�)3.s���{��_���>f����Ĺ�K����˨L5n�*X!�Sr���y���\�7����!���ͨ5�5��}��z|<ʍ��Â��E/٠��V�%����8��"�$$��{���x;8|�8�ݕ���-Z��c?�����V���K����e��\�����bh�X�b':n��{���@�C���=O�|�G[b�0�LM[�͉�u�"��缊>\��9�q��s�1��ZI������֤4\"
G��g����,�����&1-Qu��@���;�'MTy�g㗻��:�����/�k��qo� �p~�,��N�ҕ0�G�s��q����ˣa ����
�c���}���٦6��p��Ԫ춪�]k4b�"������sR+�0��c7�������}rX:��p�.ۓ�T�w����+����ml�3�CyRW��wZ{d�E���z�����RUUU7����N������j�5��ku��u����	���)|eR;�6��f�s�˅eS6���f�����
D��+`�+2�l6��-4�J˟
��fc���H�¿�i&��߳!�db���+�=Ey#����Ua`clO>O�.�)��M4+�X�*����`v�����E*�.;�����;�ئ^(���l��������5�pE����)I��pU�;n������lpne��%*�sxW�u|`�D��xh}0J��Q?~�y4"�a�m��<��e=��j31��?j��U���_�6�0C �o���~:������-�>Xai�h?� ���*�j���b:/ܻ����~]~AA���������08��Ԛ�w�ט7�1�|��ND���	���o��s��m9?h�ݔ]8��d��F�Q��4l��ND��~V�~���x+�8�>/����
�Y]	��V�֍x���Ǚ�~��,g䊗��8sN�r��F�����$:Cs��n���N�G��S�����r羱	��H�WWW�=�	����)�f�k	���Lr^Ц%U_1�F'���s[q5��P���|�O�һ[�xP�a�C��Bȵ0_#��Ȍ$^qm��S����o?�p2 ۮ^�[};�կa2m<��y�hi:�x%[��2RX+�}�`�`������e�a��/#V�be�Gk�^�	</�]����Y9�ؾ��{��;���DWc��B��E�C?��R�L	&�h��H��t='���РsE�PHP���4�`��8f����7��������[g�};��.����Lك��C�4�E�x��Q']D��^���lN7f)b@6s�Z�@��܎�/.kJi$x[�/&GR�@$����߭�#<�%ݭi�t�E�R��@��@�dĊґ�;/Q�S�����!L~�c�l�8N�z9� :"�R�-�W���I�ȷ�("��[��BBq6�A�@G���j~����~Z���-E�]��79�o��_��c
�t,
��fV�8�>�4���9��o"?�:Z5�l�������{\��?�"c��Z�I��6�ZS���R�ڃ��5�!-��O��;��T�Q�f��P��M���ڳ�拶��^P7�$H#����z�_�X�6�!c�ea"�H��A�w2QW��G )G3l݇(	�Z�X	��|��V��=��d��q��XP���gk���r�΄(�Z��?b4*�_��$�֮��U����I��-�8�#���:��N��u�=��}\4F ׬�Ѽ� ���П|���g$������/�:Uc��%���-���e�v���5Z�lJk�X'8r����^��Z;!�����N����l���42���1AQ-4�ט�\���O����d�h,����+��D��\'�#�����n���(�Rcx0l~b�1�6:׻x�0�Z&p�t�>-I����{���:^�Ȱ��JD9��5]�D�Xo���ײ��Ƽ�:b5����I��{�ܦy	��T�����������V<ؼ��$���3��rW;��ɔ��̥���R���5w�4�hDz�gGCI|�m'��[[{�b�+��22�q��?����n�O>>�Q��3��G�;5$�z�ދ:��WyZ��8�lA{�M���ɏy�w�����-]/� 'h�/�[�o^����4F$ �^Gn��`�u#�ZkS���_��Ϩ=�Qjڞ��mGVh�f�]6?�kI�N5����l�E�M�����=ڏD~%G�H��3*�ݺӤ�"�I`��'k�����GݾM[kC$�]����??�#�����ǚ%�rR}��)2���i��۫'0�r���q�ޟv���#{<������C��FC�돣�d�;��|��7P���oV�X�f�A��#Y�ץ�rD�-L�?y�PT���7F����7���R��/�x*R՜[��O�0��g9HY������*������"�9)����T����כ���BI��ͨǄ���F�'vɿ���04�m���:h#F�d��"�O)$`b�MI1��*�/L�0l]�������w=����]��*R�A����e;����Va*�@�`n�!\��%S�l o���0~�'�\ �v�n���	M6��t�U1}�қ�7OR3�S�4�v3��?a�c�y;{~�B��j{�Wn��ã��s�{H�u���PAm�_���ٽ����8�Yrd�ng��ApwJ~���fsZidܲy�)��\�E�a��dl0�4R�tE,�4ƚ�0�x�E>�>��wK*)5�-���K1w}���EҚV�k���LK~rzo��,f�[��9�Vd�ћ�☆\��G;�?$Pj���hT����R�c�z�D��a�u|����M u��=�]����?�0 $U�h��N���~�%�[KU'���L^Q��% ����+�ϯ+`��pho֚��_��fG#L�luv�sc-P�+H�Σ���g��ϫ��	
�#��4aUKWD"O��ޛ<m��3�U��	��Af���2P���Ғ��E�~��Z ����hī�xω����=/3��6X�WO_ެ�� ��Q�8�e/�F�D8�=��c�J��N��TOꆞ''(�D}��R��"��r� ��w儜�F��Z���mRC��/��t�2��T@�`��˻e�9��@N^��K�.z:�V�Fj>�6w>5x8�S�k�Ba�t��G�2FD#��Za�>�L����s-qF�sa�?H�%K�wM�6�Y������	���.-t��>=�iR�C,f��wc���wt�UO��9M�t)LR̓m3����+l/S	�<6�s��)>������{�\���Aq�_�7EAS;ܱ���WL$ztC�?���ID�+��!�+�bHV��N!�LdIp��Ǭ1j T���#ԯ���6����_.g4[��4}#i�v�ߞ=�&%+t�Aώ�I	�2N����'�[����R+���;���h�X��;�[^5���Z	�M�mMM��P�Z������� ��9 ����������Q%���|}�ǀ�c?i����lNg:�ɳ*�~��0bc��lVE�l��l �B�[�'H+_5�'�.��B�����[7�kEH����K�}�t����؝��Ȥ Qc`~�7�E?��IYy�� �ֻ�5ZaCK�t��i�`�gv�N}kkk]Ss�N���{�Zu��N�*+^5f�Msh�g�|8����M�2��_=e!�;���ɸlv�7��_��v��M�(|�6k�X�2����n/*� #���eT:k�"�wp�p�'VM�6����0�J���۵�]%2/�&�^�:E6��E��T�#�]F�{�1fi�@:����>�vU9������jqϲZ�/���<������h�qq����n��%rM�j�۪ ������88-S���C�D��j���T@��sJ�7�O���,0҇��!����zP���rр�٤{��l�ھ�T;�T�!:��/�<J��&��i��-T�r*?~�W;RoN�Z۞^`�4fd�[�N#����1H��/�g�qթ�9Ȥ� �L�&ZP�\������#����5�:�o.�&��4�$�ioQT�X��B�¤��~=\2cgO.�*^�X��I!����S������+��ܹ�y� �ޟ/4b�n(�$š�?рiL#�ؤ���RG� pQ�8���ı/"��KG76���"l �	z�g��Эq�UV��?dX3�%��
>�>�,_c�)�}�
t����D�4)2��7zN��X���?�N&��s.!�����'���
bx'oH��6,��N��G8�(�&)��q�)~4r���qO:j�PB�i�&�L_���?���. ��d5+���t�Z���o�Qٵ�����/;��ݴoo�GG7,I��L@K�S)�֫���r�>�����������V7�\�[1R�c�z�A<mS�k��~��א8��,�,P-�7p�T|Ƕ5W]k)������PΣ�ū���\)��`��Q��=(�cNZR���p����p��! ���~L2��/��M�������Z����QjUgV�@��ٟ��"q�U�U�^�ۮ�m����B�f���|��=�-����	�M}	�.x1�{O9��L����y>ZB�R��Ô��F'�B{�
Z�v�NP�s�t������_���.ȩ�� P��#>���_�]����>��ʿ�q����/Oy@��x�4��="��_	BK5p��v#��,���h��4������=�F��S�Aۿ�p�*,�������'��p��#�H%AowS>�r5B��L������z�W����gg�e 
��s{���r��Kk�����HV՞K:>�Iz\�������wYY�c.��G�������]��)&���T�9N8!��/R?�H��17tK�+�1�5�.�Oc�E�Yr-�',��Ts�����C`���nl��C�~]Sk&p��c?�Z:Dp���U!��ۇ�8H9��x�c����%i7F��d�<�ڹ�Y|�0迎D7hu���,},�@�_����%�!l(A,zz�(Tm�b ��5@��Y2�bx��4�"fMi����)�,B������`�|��ޞ���(��� z�8m�F�{̭��vOi;z�����Z�.:�z!��R#����o�������JO�s-�n0�Թ�C��}�y��9!�g8�+������dwVmuꯜ�q��jsq�qs����X2�{8@�5z��Ub8.J�!1W�B��"z=-R"+}�]Г�V���q��A QVv��ڪM�@
VH6��,*�KO�8䴳(�^
��XU�r`}4��ϫK�__��Ъ�ӿJ�:���^�p���:�
�?g.
�}��þ�~�)�_�	�V�QٰcG V�*� ���T�2�F$,�>H�h�Ӏ`v W�]��l�]�
��m@r��m��hzJm��#\�����S<g��/z��[��H������ɺ�LE_J����|�g��ƌ�A7�ھ��V�g�Nו��� �ˬ�t�WЦm�3l&�)]�h���t�3�D+}���%�gM�f�]q���j?�~�ދȣ�cX��8��w�n�PfPt�|��%�sy�:�N	����"ܻ�L�S�#pԜ��އ5�,�O�O� FH����T�[��
����	P��I����$��T���x@嚕����ӧ���z�'�Z�&��~�z0a��t@�9[�%G��Q���r���b!��D�-[Q`���'4~ld�S}_��L`��<�����[��a�W�Ŧ��Οģ/ځNh��Z�p(X|1��8s�Zx �-�A�x�ʝ1o�t�ʿ[��\C�ҩ�\� r�K�hPuu�������eĩFDB��R	N����,� �\�}O@���������"�F����O��.E3��pG��)��s��Ȅ��P��Or�\�3ۀ�g	d�[�Ag���U�hE�����R|I>�~ŵ	�߸��ٲ��7n�5���fd��X���O���D{���5\�G �klBp��Mv ���r��? ��C��(�J����)d����BP)�U�y�C 7F(�����g(ݨBN��=�ѹK{�5�7S�g6�_7��~�rp�J�f� ATj��
%7,IK����Veh�r�a��<�p����d{�d{���/�M��c��m�~ ; tE�tp�돣N[�p�u���a,ep��	��t~Z|������I1�s��������\d,�N�HZ��W6묆d&r�HhѤX�|T�/��vPk'lS�?���	l�K�"�X$P�c�%RtM�&��c�W�8�ٔA��$Z�Y%����4��	[^�]L����Ԇ��џ�vw_sQ�����y'{���^�.fp�Ŕ�"6�}�liX���j���v�+����8H]͂Y��>����ĢTiJ��	���g)6)}�B+�߿ �04-^ı,BO#I�PPP��ugUh����r�t�y�/-���h���l�ٸ������3�3ᵅ�a�d۷��h�;:�2Z}��aq<sXq��귌�?��Je�`���M�vI�B%�M./;L�mM��7`3������5~������f�͚0�g="��4ʧ\Dr[��Y�[��O�ݹ�˴�P;����_��>��RO�ٔ�bX�� �*�=��p��p|��'�k�'P���̾{ �6����ݻw�0��U�[;��{�㘋~وA܆����m���ǽl.cT�c�@��.ES��9wk��g�2K�d���J��Q�z��!,jR�_GA��;��;UJ
 
��ƈR.]��?�g��/S���A��C�#Nd�Olx v���a�h$�����_�H«(*���Ř�K���D�-L��{�b�[>D�ӝN��a=��F"���^&$���C,0�կ�����[���/��V5��T_o�����FĿ�8�� &�@��bPw[�������i��eh�A�4�N���T������}[�tS��Ѩ��x�Ъ�e!�<rؒ����E��'3����ǧ<�%�/>�p��]iz��7M�1~v{r΢���И��Ŕ\�����lU�����B#9fn���s+������tz?(���p��`�3�n^�]�Oүç��=L��?�خ!(`�=\j�I����A��)�ޚA !�X�eZȾt��1aͰb�S�ܠ�3�zI(�ԓ�仢���:5h���J�$�(H9G����HX�g�434�A�,lk�*�5|?�"��<ʬQP�y{���$��45���3Yvf X2����Z]B>��~l}��p�	J��-Κ�'P@
B$�rn�y���Y��~[;�����~���y�̃׬��rJ"gb��D�9+����KY�_(��V��ڔ�.R].�.�Z!8���ݘ��`C�S�z)���>��ٽ�%?��jn8AD���״���-]�ZX���~. *m�NS*��,za�O.��&h���W ̣������R˚�L�u��oA�Nc�� �K�M�/�O����64yL���n�.[�D2ڬ�͈���S�j� ��y<w���)��}�.������=҄$D�Rd�ԉ"߼L6����c���|!��\�費A�4�rڎ-�Ct,�ct�y �k���R!cT�|��蟶��E���XR$��@R
�#έw�.���E\#���4gbv*.z�Rc�T7홏��I�د#nt�����?h�=�,b3NN�l����c	6�׼M>������Q�	.���SK��x	�a<B�E.�Z�]s�Z���߈��� 1��֐�D�=S������T����V2Zf����H[���ZE��\�"ԕ�F\{��}�E�-���е�_o�����N������|�����B�T�����Z��KS���<�?�3���%K�V�A���+z�Ϥ�q.Q��':��?�ُ�=�׿��84>ZA�.&�
��Lw�!\=�3�=��'Xc�$AЙ�%����1�ָ����^���7.w�d���C�),��I.qʐ����{߯�c ��p��ҝ dj|�a�� ��B����Ʒ#��~��}gy�oqg7�C�ڌa�m͡�ÁB^y����dv�;��i4�5��]�\~!��Q����<p]žEc��>���P���c৞���4�8��̸�-����L2����f�;t+󉦔��F��l�dK����,�ݡ�c�pg�E�iR���#T�/��ۑ���fQ�)�߈g�����^6�3����!�bE~�&��ş��X�ؼOkג?�����73>�����
Z���u��{�旆!�������oP�ܦ�j��0���|)l��S'`S�P��?�S_s�p��J���9����d[�T��,�Y�Е�{�QW����<�G\��,4�i8l�A��͢��Tm4�C��3�P�$���g�CE28}��З}�tZ,�L_%�~�Qټ��]�F�cv"T_�:
5�օ٬0j��S��m( ���1���61���2�)�৮@>|�	X�[51��;XSwy�QG��\a�u�?ſà���Gg��& �f�Z�% �Sg	�`B������9Ȇ�Ш�X���7��x�d�	�n���!��o&�P.��.�ڮ���e��
��K���G�	�~V��}2*c�UC|Z��Y�����B��$��F�5 ����7x�jEct��݀�l�U$]��{���"]5�~���B]#4��acN:V��OZ֊L���ts�Fi����5���	z8�N���4��2RLD����1�u��~�����{��f���,;w������Y.��aX���bE��������F+��n]�/5�����>y�[G�z�J��f�!6/|5iv���h��Ȇhሃ�;4�#�}�������������Fb��%;��DI9��,��ڧ��v��]�,�z�)s�97 2����DLQ�dKl�U��9!HoI��ܓ��J�.����E��ܜ�[���T��{�E9�c�����W��k&�/�CշEA���=�%W����_.I�s%��~�7 \�:x\�|d�U���W����c�ey����'K�._����B���/b�����E�^O�F���"ԗ�"�� ������>��h��
]. ��ؕX�H�9�E~)z�ցb��0��&�LŹ����_2����\y*������W��������JQ��dpvr��S$�,I!���r��띾�h�&`D���&�;�i�J3����F2jcû;��Žėc	�>g�c�ZZ9��O�Ζ���5Ł(���T�|����`B�`*9�D��7
h�������1�/I�e��4(�$b2�6�k�]���:�y��@wN���B�f�ϒ�>�(a���>W�=��x����R�A�{8�3�����/�C~�4:
�8�^ӈ���}��:c3����>�"�-��ZhKЉ8+r=fj3b C3}�_����b��c�ae�Q'w�2�BefJGcP�c�m��Pz�q.t��`�%׼c_;��?�]���q���{"�wHE3�VO~(�|3�~�j����.���g�x�*��*,G7���3��q	/�Z�:� �uh9fA�Yb����@*S>F���>:<�i�X�I�-���W�����/��>׸Ys�S��7�7Ug@����h�SrJ���袅����!���>�&��M(�7>����l�^�H3z��sj��g������;��,4_p�DW'g��;Vfl�t��|_[.%�m?/d�?���8J7Tor=8@:�2(~�(�R�W� u(	���W	�Ǯ����`n\<p��B�
�-��~[㪙��s�`���]o��$7��O�v�G�<;h0��^���S�_)1���>�u����&�+��e,�R4�:�Eȓ��W
��O��$���̠,D$x|3~�~+�/ ���ac��$R.�:�
p�7�ǲn*�:�����i4Zjb��k��rJ�:�>o��R�U��hdl"�P� h= 5�k_�f��A�6TJ��	��R:4�s��ZvO���M����K��5��O��3`�X�y�y��	��I9"^�E�Կ��x�g��@,(L:��,*�n��s�$���O��$ʓ/��
���2O���=S=�BmBr�a�!Q�?�n	�٨h���������<(�x�~G��0)a���bXu1��p���"g���R '��������E#����=���**aE��O�����~6ό���׀�u&�=�и�<`�գ1����_;�)Bc�}���Э�~W�)I�O�a�,5*�*,1�1��a���_��'�I!N�Ms�f���ޙO�;v�-�p�?SL � t���U��H����\�e'O��%�H�E7��#E��H#�+�>��ܿ�cH�j4��cȴ1(�
�°�t�)z��;P@5=�H�?0y�$b>�)&�S 29��`t��`K�T�bqhss�}���F����|{N��p��r��L����L��f�:;��sB���u�����,�E����+���z,5Z�m�Q7��\��}�e�B&�0'���p��-N&�(�l����?&��āl<Q���5��c����i��w*��iSrf�wMxI��UN���W>�s��� .�"
O�d8w��er+����rJ�R)�����1¶I>�D�8�<X���:�_5IIո@����1sS|I;6�RDq�: )�,�3m�p9'x14�#���ƑOY'��!�9t�5z��5"F�!�����;����c�9M�wt�����8F��;Y6~����J9� �BY7t�+����lY�m^8�p�,��E��X�d����x�u[4�7�8�
h���"���� �{��w,,�;���r#�S61$*c��IP�

��И��q%��Q�$���`__��X��a
�M�ad&$��ᑃUd4�c��9��A���{I�;�����ѐ��$+��@������v�.����&?đ0�@�e= kj_m�����xX"t��$���bݑ^�"��������@�+%�Z�/�?mѨ�֝�&;u⡦�͔�{�=9CE ��
�Ñ�K�@�@ɻn��X��R�t4��L�zG`�ba��D�S��w!���^vݤcoBW�(3tX������Rʬ���Î�^���JGޞ<Q��s��e�9��$1I���PRTU�{d�����7�[�˷�y?Փ�|�I�XF�޹j\m!H1x_8R����&��N4��U�"`�>%�Et4X&��G����{�w[���}z�
k{]�[�{�0^/��u�[-L~B�:1�;m�\�IkO��^��@s�"�p=�*@u��'��M�˙F���C��d\�]L7	qp�}|�{��1/��'�G�CtF�ߪ�L-w�}���l��%���^J^�ey��z,N\\��|N�i�WT��Β;����B�T�e���k
���!"�P	r��vbV�yu�_�]h�%��K�m�f�����Lx\xZZR}m63`|�J-9�r�N����l�{^�9:��U����i©�'�<�c��"i�<�,`�oѦ��ﲗ�y���Nw�Hɾ�9:��}ΊH��p�H6&��54ۦ�_9"����+����t�l�x�ĭ9pp�J{�}�p^�{���J_2������/P÷�
������ ���5�!s�:!��l��'�L6s8�*=bʬh(��ur)��$O/�H[z���C�>X+�Q��gX?�E�z�^櫳���`:�38�(�r ���T4����?�P4���3a�!�K�e_��m��2ƅ\Q`{����wq#�o�������T���w���WS��(�h�QqoT�@K(1J ��&Fp���`8I[�I;i�8
L�K��~ʀj��ݻ�\WJ|�V�/����}����K� �"oh�SH����_%�Ţ�B�v����w��7��c��6�ׯ�c�F��۝"01�b���"���B���Ξ������.txoj\3��ãz�O�hB���qYG���{��(��d__�$�����ih�F�l60���U�8׸�F�!/N�PM�����G����@�o�2�<	=ᾙt�6|�8G��z8�v5&���(�ިq�⥠���N߹�&�&J����:;!����Q[7�)���(��y��

&������A��]�3@W�Og0����
���J�-$v�B3~b�2b�|��i�N����,j��ǩ�����w��0����&��L^$;��
ੑr��D���dQ�S�+ާzUu��S^�?��]�@?�Ky��*���4H�L�8�	f8[jp�B�/~������.>���b����|"���q�.�5{������^�'��	���m`��jz=���-�x�*z���۟gd?q,��#�X��(|$�p0U?��-�g���E{����er1h�?%*�H�?B�-�GS����]Q�/_�GU܆nA*����;W���Ls���!$���C9ڱ_������"O�U�H�& �?�=�_
���\�zd�A�)��㗝	��7Oz�:��׍��3�vjJ�w�z���ئ?F��kl504�e��{�W�sK%AӉ�F�ŝ��w���ûζ.�����D6[�!C)�^�1"S���L�#�`���hm�荛�Z
1bv38��B��>n�}�(q�TQaoc�+t'<��ߣy������/����:텒�Tg)h޽�p�� w�=�K��7ۗk8e�@J�"�$,�&���=�u�{�tc�7fzG?���ֱ��j٠�w���j{�Y�kO����%8*w����<GR�n��hc�n���T�/�W�^U�A�h·3�*T �TK����W?��J5���D��� _�E�{�'8v����	��&���dI9:'��As���^���(�Sm��]q	H�#�]����!�
��_���ip�B���ÝUA�v��,��~$��aa������9����_8����/ۧ�������_?�o:�|���ၽ��2?8�C����	�}x�i:[��y���0;�$��'���GSߥ�Ε�����/�w����<C)�g�*Vy�����c�gy��ˢ��dgUSc9� dB�2�۫��R�ˀ?��(E����m�V�st�uZڝ�P4������_X�N��(z�MY�sM� ]�,����$���$�����:{;�UC؞�s��e�Q)$��.�8K�7
��=47Ϡ�憊t��|��E�=?�����KZ*�=	�ޠ�s�:��l1���R����bj��T�>��C����ZJ!����]o���(��"�_�|B�ك�����G!�+f@T9�l����A��� C"��N@���9x� ����l,�����J�0��������$������w������H�{l�,�e%�L꽯8LR__ߨʈ�̚\a`9�Z���c<DBkk~����=Ѓ��s�%�=��=��M�U$�W��/�^���-��2�v��u�)�)��?�Ru^"�Ǭ'��#[�:;M]�Z��kh��������7������Z9��ٗ�De����N�'x�*��^�~a�����f~|V�+��řw]������Sg�ST�vZͬA�&әq�*�%��T�vxx�a�֏~���D���v�S�`�ꂆ=��6���_?�����W����H�h�Ba�����!���4{"ۊ�i�4~J��+en2��Ěf͋>�S3�� �j����iF�	�hP�H��-j�oZ2���1\#���N�M��l�]X���$̘���u��7����&o��]��n�^f\(~q��֘?�����ؚ��������)�UiQJ2Qq{O�0'C_�X�NO8j��1����A!
O0��A[Z�\Z͔`V�>Kj�/��(�E��bȖ����MD�S���K�Ey���b���VE~v1q���歳`�*w�oZ��Y��߼m�Pv�P"_�x�n/j�=N+�5����ϟ༸q�Gc��pt�z^�lR�,:99i����tdk'l?AA���Q{��wТ� �F�.��>t��^Ԅ0#��h�I�`���r��7F2���G����[MM\����#Y�d���|p�4t:�5P[8%�'�P&U�vC[�B�N�)&o|��&&&B�@��GB�<��Y��;�iM'$��,bo���MXCa�t�!X���0
WuA��s|L�G��Ci���^8v���Q����4���5�i�`/2���	<��SE;t�C��D�@����4�U=l��z��Аe!)Ŕ�"C���P��@��s~]M8Z��qw���o$���0a��go�׏#�s~��N$��"N�b�uH�x��CӦ�/�F�j�У-EEE���<�U��ΉY�R��;��c�����
߉���_OXoŻ��(~j��5#x���;CΜ��;¢P�9ă�2����_P��X]]���}�뇡V�o���D܍ T��|�����ih��0-��
�6ι@7��5�!Q�#5�~x���w�l��y�꟏����ە����(__��������j�%q�y,4��nTO(Yh��o���/�㷭���f��{�>ڛ*}��l^↝�h1�|���O�K_��]#))R�Ss�����}7O��,�j�/[/6p�P1;w�s�1⛶Q;��lS6޵0�?�}o`p�>�F�����N��88^>�-�[Oh��+)�k,��MD�ׇ�I�S
`�,�T��nJ��+��|yMM��DJ��j����� J������ǀ��� �O7Wr��!�8�69C�?ws��~�����&�Uό����3�/�Mĕ �i2�m�p�z��2�3�A�J�F
+�B��D)�ǿgS�e!���$�L���Ϧ�{���R�d�7p�Q��LM1M�]�:���k��#����[�܉��V��K/(�ry��`V�F�l����ki�Έ� և�D�zf��!��GM���}�!��'/��K�<�˚�A=�q�i��ё�H�:���h�14�7?m�,2/�_Z"W8���X4Λ��Ѥ�ݺ,�;�u���$��=U�L���N����7�I���V���o��af�,*H��m��q�\��ntM)c��#˕�L���w�gk�J9"�p���g�m���$Hީ�y6�  e��W^_��ӆ���*R/o�7���LS�J队���T��_�A���*�|�>e��yۗ�cT�X�
�f�o]�N��N>V֮��˗G��Iզр������(u�2*i�w�|
�R��s���P2
�f���̑Y�8��KY֛�
;}ӫ���_u%r�H#v7�-|��1���V�1��T���3�&S����-��~����[4o�zz�n�rwwO�����ո0�Omqx����~�Z;��:�Ȃϻ�ƅ�;�����I���[���5�1�R{<�9���~¬�0,<q�{� ���jd��W"F��t�2�z���^���7�*AF�k��zt赙	5I�� 
�M��'-,|h���,B�\iԱ��nuR#�͂Ỵ�-�#��8
Mu�'?�:kk?Yr���P>;�I��U��� ���a��Io>G�ڙW�5��՜�6� �N�k�h,��W�m������	xإ�2���7%��D�+a�"Qd/�;�x�3��O�c�7�O�GAՐWP��"���ق_�/�^�)�g^��!�OL4ϯ�Ȟ8��%ti�"�t�c�f��&mn�Es{�b� bK<S=� IG��jהOm֗�KZS�20���<{�:�h��(R�~��1�N.f<u=��b���)�W���_mFpݩk{��B���ua�~Gm?��n��K�t��A�I�������림j��&8�"8R�;�[�n_�L*ICS�%��~?<|������0���6���R:���qN�Hd��`�� �}�y�Gt7������D,5Y�8(�2�_[�B�W3�8���}8��|��#h�Y g����`d:KA���p��N˦��0�ε�~�6��jm1ֲ)�[k.�%Ś!�fJ��3c���tC�FFF��m� ���B�N��Rf?rd��TG����)�����M�D�H�.�s����A�qXx�Z"��ن��Q�w�ɐ~4�`�G�n�ӑ��1�~�<��Z9�|��37B���b@(;�Y��x��;������mL&��k]U��\�媦�F��s�20�����g-N�x����6�;�p��`���D���D�n������L�h6[7�Ά3�l��q>8�g�c*��J��ۚw�$>)���?������}�"�h�O��0�ą�
��N�cy�L�ΕH�� ���?@+K�|c�|�2<A���Z�G�тn�ZKu|�ds��E$�U�a��8]C+�2���p�����5���������E�sqX���7��!5��g%�{>|�.���#<��A��*-vzEO%~n|��w��i%��&���T�:�'_�A#5
Ŷ�{�����m�[.���������{�y A;�׃4�V��`�0�C�m-u��z1&rf*v�|k4?�zGcp��]����@�4��zg�\�������6�{DN�v,I�^Ki�aV�G�Ld������S^�� 5Qvt�o���+4%}=f�K�g�������7�൪p{v�%�瞱Ǭq�8�&���\o�UR����~���QƗe�[f�����RQJۺ	��S�a�JŏVIۯo4�$�)[vg����6?�Z�s�y�޿}L�!k:����o,]Vg�����<���q��ӬϰDlm~�m�J�Xm)��Q"���+w��9x�Q2��xskk/�壍huv�t0X��R�[
�>����-�a7�Q��ϴ#�h�� �k|�M�WSS�WǽX���'%���_&�.^��+���kk���>���g�d�~�鹸�FKٔ{�8�[�L��l{���47����5�yB���V�ꟗ���D�;�$t���/n7�+����9xvѩl��(�����2+��%L�џ�J�K�A�*�ڤ�_��6���=����[O�b�&��ws�m���"��M�� ��#��n	�d�:2~fN]�фh	��P���p!����j\B)���!��B���9]������O�ɚ-o����_go�Ā�	H�J�P�>I�/�q4�Q���!����Ё���ul�FU)jس��q~#�[��]�'���<mV|a��/����eW4z5���(�n٧V��T��ߴ��^�i�/�^�EG]��G���޹N�~�b�K���M�5��n�o ��7�_Mp�E$�6�c!ͅ][�n���JW��^�P�B.@9���e\� �A�6��Z�K�x���b�MsGqx�:���k����ƒ��h��
n_��`���qr�PwL�m��R�Cy
�tJS�"�ym7?r{d�t�ٻ.-@�:�����������,�7B���$��9�u����X�X�Jyn,�ߚ�1|������5#N������5KLϥ�e'�mb�t��^��Sm�۰�[���[���]�����U/�BSc<*߄��T����om�s��\dd��D�����R��=m��#�q�Z�����n+�����e�L�_�Q����dk�b��+�-����H��X�ۙ2�����ȭ�yU%����t��Qz��*��],� ?ou���^���Bn]��1h9��T��D����I׆��wC�Dlv������s��sن/J��0�fz�I�=��Ԫ��G���(TH1��)Zh#kt�R�`�4� qxtѩ���#��2��=�E<���s� `tE�>	���fӞ�y��'�΄\z�&��Z~t�+�ўX�|Q�/��l��D_Vh��X�S�i<;��l���l]��97?P���r:�C�_j@�Ve��ȅ��o��ثu���R�ᯚ6~�6=�җޫT�U��af8�����~_!.n� ѤN�S���w�8�y�m=� �rۮ�YS��:W� ��-��F�$��D�]��7N"n������`��M,�Y6Wۻ�Ԣ���sEI3����oztˆ��ԕ@����g��6��h�>�n\BiZ@}|���
����vvBs��w�#�`B�v� 4-���7%Ƣ`�����{,��V�{��rW��}2<@$o����:Ԁ�����"X���z���\�CYF�+TI:�Դ��O�����G�M�2��u8�v�|j�H��!���?�d��}�O0Fl����=:�G�}�C�){���ѐa�,MJ�Q����2�v��P=����R�����ϗ"}�L������!4��`oME�S�a�[��y*��G긮}.Fh���^桇��&���W�աz:;���K|9���#��1�k����Ҥl�>K���=����j'n���|q�/�bX�ܛ�l�QQ�۷/������tR����1�+��ܪ"��r󡎀��|�����*��٧��	�I�k=�V:��!���]p�kN a��$<�-:��r��#R(e-�gI�
�AIiiO��qO��"�:���x�!߸�ܱmm�'�˔F0�yw+(����~fy������[kZ���n�5�_:��]<<�i���哪L��.�v���\�����[*&Ĕ[���{g�An��Tp?A��W4�g�Ζ0r̋\J\B�����|���7���7����_n���O^�Z��\�L�.J
3��N���aI�;!0in�Va���{��&�����K(�0gd4��|�h:��k�K@�O�d�m��J���h����ʎ�3�l��ZӃ��WV��P5��xئ@ڙ��*v\��gN�g��1 x&�F��'��aE�Vyj�{���>5%�3�vٻ����{`�-N�)d���}꣬m]��P�i�V��<p;�񿴟|������b��usrz�3'�զZ�xH���&�ێ����V����H�����V6�w��x���S��S{j�?�ȼ�_�}Ɣ{��a��yf�M:d)v-:ￛx�Q���*Pp#J��������Q!��V���w��9O�4ϖ���1�>D�S/�����]�������H�%�>]���b��J�[Y�ۥ�sN1�����ݨ�/&0L�sy����/�^�	����*����֪}t�5�]㯉��ޱ��Ah\���ݶf+�3'�bemYEr�� ci�^tdѕ7l0D;o��vi��w��&�T��t!�p5k�K$�د���4ߕ�Ȇ��x�/*���/�����!sDg���~|���ƍ�/f�	a��^j��SiD�J��p+�^�		W��(��Pk��Ly���+[`#{6I���%U�r���R�/o�%vQ��Z/lv1��Q�`�Qv�J�hsrNj�Ϟ2�ц����y�W�c�և2,�K�;F+nʔ{�2J

��3�Hc	�R��$G�BF�n��ϓ	�AO?��.��N\ӶT�y"z?a�м���ߊo�@������~m��a&�b�����[+t�:����@���8�3�����@�#����{8��n�TJ��XbxR���?!�+nIl��1�����wG5�@��uTT��4P_��Q��r~�	�qq[����F4��Q\��ص���ke�������Ҳ!��d�6�:���1kݶu�X1�1����m�v�X��(Q��\U�p���������+Q3���y[�[V�>^HLז�.͛���֚�r�<E�F���i�=v�B|�5��k"���w�����L���Y�ؒ�z��3�{ ^��.��k(S�9O����6�S�([��,�`�]��wN�%����H>�?����|�r����6�L�R4��_h�Ҁ�DG����ǖ���C/�B��j���!���󹓓�r��/&���g�V��e@Ơ\۝�߭�{��Q���=�� �
fo�6��VL�)����K
�WU�-�d���Z��z짶���A'�-���im�#N�h��ݛl�49�`[�����0��=i2
���8z�pk����"�U%�#�d��������5��b�3�@9�V���Bm���N�e���Ύ�'ۣ�1-��=�����l��	�5�;�$5��=���c\�BSH;2�v�1&D-sz�:!Y�]�m�+)ϡ��O���ʚ�w�R����'S�U���~�sh#oߠ6�;7`����ߗ2ͤ<^8����t��H�lL��M�=�����+g���({{�ܱ�k}��3��!ʹ�΁k5�~a4}��!��₭�	d�^�_��:ў�n�$���!j�Y��#��8W��/y=��HKK;��%R�KC�]s��R��C�\�.��9�ݢ���te|/��J���=���8[ xff���X1
7_X�EL:kQ�]#$xS`�l[j�M������*べ��u�������ܱ����;&���lgV���**'C�S�_�O{~�@}eP�3QU]}6�]��v�����ѽ�I��]Z�<�'ݨ<@�`tD��KJ],�̩EO��mʕ_H�D��1U��?NG�hM]�ϱ��\�iK�Z�k��ы�ł�'�W7Co���:�`O�Ng0vvu���Zym��^�;;9U:�d�.V}�H��������d�%Q�����/�ɚX/��Y��8�W{�@�s]�K��5�8��!z���r!]	^w򍍤�Wv����O�a�������<�$�8\�=66�r�Ն�iwW`�fi��v�^�/�����iY�Js�X[g�8�������S����j�Vs�������������h(�^�Q@g/oР���e��� }=��X���й�a=���p-K�����l�z�F)��T�4?ĲdX��O��<k�r�J��>�7����o�=���0���P������J��ö�]j��?C�lM�̩�6��u�PҚR딗��d�n�91���
��eϮ���t-��?R3�S��4����G�YTm8c�N�[�)J�ν������#U�uuuМ|�guqE����b$�-	4����9�jJ2V��Crn���f4+6��>��GP`jjj��õU��?�_�h�>��㙪��k�F���p9�:�����_�ɘ���P�Q�Z��yP���N�S�hjc�ۋM^��t����맇��ˋ�/�,��c��y�,���s6��lv�9����tS�����
`e�]��(]�P����QQlH��� �U/}6ܘ�h��R�9mĘ�d��f�$���4�[i_�]_��)�tw��)��������/x%�߅��T*_O�b�V���}J�س�j@9��1�����#�2��μ��sԎ�l��4��TR �~j5hju�d���|��O4�\`�4���W����0P333#��J���eftv꽯7a�C�&4������@�QhR�6Bj2�~R�i%.&����m�p��N[��[���.���u���� p��sSRO��	`Z]�������tG�?i�����>H&zTKxn���p6(!o�_u��d���:��3���5~ȕ���P��d�i �2d�k8�~Q\]/;���iy��D��_]]��g����� ��ۗ������f���<q8��?�j^'{wgN}}#T���	4s�sV_�\�{Rô$�4Q��{���~�q=�mJ(QU��-���7>�p�a�jUԅ�Zf9=j\؟^ϻ�sK�Q�"f�\k�[���_����ƍV�L������J]G.q(ΰc�^��b�@��D�|�׹\�ܭlI剉�@!��a���gΜ��033�sT�*�� ~/�2�ATWww��pCn.�����yc�����������Y:��glH ��+*)�?{v���,�R,���L&���H�3�b�^l����zzzofX-X�̡�4��dB��v<3���(�>=5777��i��-X��ǂ�%��� �0�2c0|�~Sߓ�t����O�r����ϓ/�Fd��K�`�c��s���z@B?��z����($�A��x#G��nF�:d.� �b��J����V<��Hv&����lgCj�i`���Q˻�űB�m�#Ma��r�TjKu�\�ˍ^��s�$+�Z�A�	��ŕ�/,��1�*��xM9M��G�d��d�A�W,�5�M*��þt������8�\�З'�ي�;׶�|�������(��� tv��ܼ�����&-��?��?5��LWW��/eۮ��/�er�G�:��:- %��y/�<Ew?��j�R����ِWZZ����K��}����ǳGmI�VZ[[�Ԋ~����^=�?��Q'���={����q��{��@����su�N�]����h�$������{N�-��'R����[��ͱ'��q��<Q����Q�B���A��%����n%u��z����͹�v���\~�&ό��o���j���gS`)-��"��	�����9b>�
�OX/�Rh�UBq���3}��J'�����0���'�*  ����^��b/rC���;��/n�L��S�cf`=��Ҍ�-�M�nħ֦�~�c���O��Q }�����H����e(��q	�x��E"��R�|�
᭫���:���߫s�\���y9������(�]��*�S�+=�9�N��瀱��������a�I��{�6~�Ħ�-��Qi���� ��&8���db���p�唕�?~� =ǹ�����Z+/$�O}ȳOT�� yDvnI�Q�X���Yu
f�]���V�5^A5@�u�Β��-3Ù'��@� q�T��g";;� `���v��b��Uy�����.�H,7�ua�[�4��ұ�þ�$��ϋ�a`��P����j�q���[
=#�L��3YJ5Ⱦ(����o���{�x���}�Q��;�Z�K������/ġV�ΥБ���phMΞ�q4�ąTbk����ƛZ�M�� p� ���wOO�l|��ZM�B��!�%ڷ�=�Ll~���5 ��� ��3h߸�֗�h<� ����鹨Cj�t}/zf���̀t4#~���P�!UB�X��6	��K����=���&��,�v���-;�e	�r
��uF�e����`�|���o�O�����P�9�6�W�RI��Q_�m���C�:
�������2ٶ��Z�U��S��\SR��#<L�EJ��y�yM�蟹�}��M�{�4i�2�>�|V4��].�B�y˜[e����"t�q�_W|ȅ!u�U���8��Lmm%55)�_���������Q�D^ޟK��T!���8Y5�����@6����
=���g'�{W57��5U��vil|{��-����/~ �&��⁢Ǐ_��>��T=�����Z"����5��#��>���o�1�J�[Q���|7n��>N�_�	�f�]�Zm��� .�'�$`����!X�Q ���n��5���X�t�z4T?"�T���,��2$��K@g^������h
���X ���r����a�aLH�e��АÓ��p�r�8�rnccc�u$Z9��$�Ӕu؄7� vf``xY+����a��[?��ɇ�V��� `�$a��ڀ�{({�b�����UFɔ����І��Ng����������[)�p;"����ҷkg���|�slM���-�!�a]e��>>�@!��mU�^���0�+�Qs h`����X�J<��c�0�}�]^.@���tfSvi��j���/�Å�[7u�;�GB�WM^@ɿ��Z)8<�7�r�5��8�����,s5��ҷ��,���M�@����;�œt�:���Ҳ�����pN�tT&�}�~mt�(X?[������j�¤k��M���#����+�^~�F\i�]eGj���ߙ�,j�8�|ȍ �իW������d_(q��xω�@���F�~]�^L��������{MK���><-�&�4��4��K�苖٢QQ8���%�cOJ0C��g�12r58����텇��,�pa�o#��絛lJ"�n�>�tF� ����JS>��O�@�2Ny#=�׮#�!�y2eM~�(�,*(�x�?�uU+�=\�������Fȥ;8�{�ahO�'��痖,""�O��Q���'�T �E����h@�^����p5��H&�TV�q�r���\MG�y4w��V�R[�=�b��a�I����qC�U������lH���}�|!�뒂Z�t�6�Ԑ�U�_̢cZ� �����S;�n��.����j�CVҚ'"̊�1RHT�b��죄����Zs��س�I:�R�%U�%�E��섄���)p�;v���g�H��������2��Ѵ�Q��� ߛHUn����@|��(��6�C�Er�^/_uQ`C�7��Y&0p�_��p���P��*dR���u���!>�^������	��k�,�^yM0QΦ��RCbЩۉ:?��6g�Nܱ��򍃜��_�Ϭ���[�93lcE���%^����	�܊�S�ڗ���Ԓ��#-�dX.�j��ȡ8״M�Pj�{��� 9����YYZ:��t����5m���7�&B�B���ˠګ���y�ܚ���*~1�O���j�`*�F��Onz�,sZ
�%A9V�6�,�E�+~��#`�r�6a){�������^,���
(K���f�~���. \���,��ڼUUgۚW8O�z�?���X$�c�B7?~� >��e�5Q�驏yB��Df��I�<�KĎC^��.n�C[�U�xC���g��l�`϶����a��{k@t�	Fxxd��_��h���u�
v���rHc(��z��̣���4����Vm��E�մR�B�02�s
֣�߰��C�lWn�\�S���#H��s�{�>�M6(�B Y8�;�y�>e#�>}��l�(�v��	`�g�%1�y�Kp�T����<Û#'���A���a�!�7~M���o�zj`mt������+t�����X/̞�x��%_Dkjqkj=�y�IJ�Λ�+ŭ���u^�5Slp��mwww�����{�](��G�wG5�m_QP�*
*M�WA�tD)�"�z��Wi��@��Co�ti�w�Z���x�{���;#��:��{���<g��.�H��7���Ձ�'�㇛^G&v�G�z��mV�u���X�A�C>sraX$����f��"*Ɍ/@N�8+����3i�Z}� w�j����g�m����$��;�Ȋ�i�	���˂��l��:�y����0S5��ͅ�Ψx�D��-99y ���M/.5
&H+mDx���y �@^?J � H�p��٩��1�tM5�9�����>�/W\�0���t�ޣ���vu j����>��8$K���A�%�DtC=�&�>Ѡ�?ծ?d=�o��W<_	�P�5!� /����̄�����Q�A� ��ҶṺ�����k�U%L�=$�g1��؏>ܨu���M�}��@�y��
Xxtm#�s=�H�!���&~�r1��=mξ�)S�ֺ��H��a����/�dn*����x����GL6޲X&��ȪC�f��j6p�����FjD�ڜ'�t��S��JJ��O�`_i�kul���5\u&{u���Qo����1Rg�0mVO�� F�sO��6��WQ�jW�^c[(Y�6˱4!����̺�}���WkNM(�
^���<x� �q�$1`��@�;��d��8�.E��;[���t��7:��*��'��#vD+�XEE���u���o�ݲ]��H���'%x�:$�p�m�06��gYh�o����y�Ԫ��Ґ��(]�΄�.gܖ;������ׅ��zd����]�!�`hr2����}˒0X����cڠ>(����U������0������8����%%gr7'CT�� D�:�M`�n���B���W%>��SM�Z��"�[8����Ĭ�ri�ٴo�����^�a�}Խ�*лt�`ƕ���m.:S@��(>*�D!�/�\��ƻ��TB�oo\��^���/�*��Č�2��´_0�����#��&�rUm�r=�X�mOZ��.�a�G���:��Q��Z��獰����6��Q�d�鱩��:��&�Ǐ���WH�~�-�r�z��H�%�&g��5����Tݒ�����*��c����缐z܀Mn����r�@@xʗ�d��2<.r��9˱������mf�!�Ɂx��]��͈s�9�0�]1��"� d0aL�k
&���J��(�U�H `����K���g�� 0j��jmm��~9��t�]�~���a3~&0p�N���o#��P/��H|��4��O��tu�,G�X�����R�PC��i1��p��4"�3��$%�CC,��ׯ�]�s��������C���-�PC��Nn�#ڻ��%�Y��7�.�M��:A���sċ-�>}�/���T_�u���k"�C�<�g\o������ram��5��C�/����o�Ex�nkhh�|�:02�[:ܠ����uh1Wo�b��j�� ׬1bn� p�F �B)h.T�܉�xA�@@,aA?2�Nw�5�%���^�>N�`����8Ghh�j�� ��!�]`�(S�3S9���w�׏����fq�R"�)�:�_	##o?�ց��mYI�1��Lr���0ĬH����	+]��0���O�H�&�~���H��ӻ�}��y!�����@W�������ۿ�ۜk����ȑ����yyK�,�U�;�Z�2��/d�)�$#0���@�X��Je^lF�d���� ��z�.� p,-��D�����e����Y$�6 ހ��w'��A����ېSYY�05LE/����u�.��_�|�~�������0)�N2����RB�"���Xw1q�Sօ��=i��K�3O�JlQ�S��)��-셓���3Ņ2#�;�=@~�R�2��{�qVL}Οh�8��ɿlW���h\�5���["��=x���zl|�9%$56:��d�@�Y�	bl��� y�Z��1����>�[q�����~~���#U�+Z�K�:�:B���TI_���1��rRz� �d<,"�#��ҟ�8A���x� ��J��m�	�� ��k6�2V����D%6!�?p��8�����G4�-]1gC]q��0Pޠ���Kݵ�f-���0�a^2� ��5��v�H�
��Z�n���g�֎�)���/W�h�n#� A:�Q�7���p%wO��i�i��W�e�'��w	s������^#�������hL9`��W�>a�!%~n���_���N���'���k_�C� �P��[G{I������`OU���� ����0�W�*�v�Oy�m�.�.�����$�����A�փ���t�m��ʣ+Cx�%���H�M����Y;���Y{o��������?�����jJ-��U���M)�^��,�n����܄<��FH@��������|�Zr����?�����1�Cx\0l��[� ߸Tݯ�������U!����kxnz-�%V)'V5/�)k��;X�� �ѵ���~�Bj�h�5�F�D�'AE./[g��&�5��@ٍH���D��{N{��`�����"Z�Z�i���h>��	��ar��������f�Cg��Cɉ4�r6D�S.��������i�H�'�o��q�B�D���^����1=;��`,Zjb��(P1��Δ
��w���A�*�����)�i�}O!@mJj�uU�3�у ���O ]]�d�:ұ�~_��Q��Чť%!�#)o�hE�ħ���M�D*�M)����o�~�z��y�P7ˮ�a-�ccЕ����P:|u�B�/~'��|��ˉ.��a�6E�r��::��Smdr��N��ۻ$��?b\p���Kx�LY���H��}Eհ��gFq��9�t�H�È�U��>�C�90�P�&���ob�`�cE�����r������4S�����c�*���l������#�=�=���n]Ā�JO�<���h;b^K4��M��n���E�~�JK�;rr�[bd��Z�I*�:�@59s�iH04���#�_�?t
�����_E_9F��q^W�����ǫF=bcW�Фl��/(Z[/��Z?��Xf^��Dc�g�Z�l�ix��3��L97_^Y[R���٨h<�����SO=���C��[�~WG`��<����6K��tP%ǁ�ʻ�⦧���f)�:&�p�%�1'��� ���А@y�3( 4��1qj�~�\�6kP\�¼c�\���@^A���̃�B�x�I`XbI|Z1�ڴsaK�ƭ�#F�;�7� ���{�_�A�:zR�	�ql Sn��+[�%F��c)��,ĉ�"�I��ib�5�QHz@�^�����O����Ǹ�h��l�=�&�|#�#ZQm��a?�b���ǽ[���h����[f (t�2�P���`��Ʋ�:jH�6�-���?�T�/Xr�9:�51������ˤzڂ7-@���K�䮑,p���"ZP_1�5L~qt�v�~�`��A�ݘ�U0�bg��g��@��}(AQ6 �uz���x�ϩ�)�leK$��^.'��h������%��Ռ��1C	����X�	4����I�B�=�߯/tm�"���P6��wy�Y��բ�D��5H�JLLLZ�o���hUa���&�
��3���Đ�W�o�h�+�G����n��)-8���@��-��7T���y Y_h��w�{��~O�QdpB��S�+Y�آ^??���h6�p�D*]J ~�Do��CgѠM�8µ�����!�=��ߠ����f�x���e{�"$���צ�ѷ��S��r�_Lv"��%�+�7;�oh�m��t�xc�ֽo� ���� |�����@6�K*����hi��m<๧�?���^I�^�j�����v'Hfm���D����Nfff��(�/ο�@`-hN�_�N��F�(�&�/W��p^E1�pQVL>��DT�� R;O)�P�x��
A��'��BD D�O��g+�v��DFxu�"+�?EG���C�4~���BXa!�e*�C{�TU_���&^i,v}�8Bg�4"�U~�<�ژ�J}OKpWB�<&il�8�h8�ڮȚ��jNd�������U�~��1E�3a&$F�"᪭���19�"M�3��	3���+.��ц���옗v	�c3�*<��U�����{���#�jL��%�%�C6�����6��j��+D�2a�}T#-�]-dj1M����Y|�����!�zkfڄlҩ�����bNB����Iָ.��Z��ۮ��<����d�]�1�/��ȯn�C����6���kʋ��|�\RNlQ>�H��W���0�B$����8I�O�w=:�!C���S��#0�j����w<!vހ/��ob/zxgb6��<��L4=a0;�8��|뢙�7h�ǖv�þ~��sO,*_�l`�ZiMI>C�^V<Zb�HI	�{J���uR�o��� lJ��bTN��������C��YZB
/��'L��o��� (K�1Q����'|FE)�|38l8PHj|x�8$.Ņ1~�H�#��x_��o��7����n?�oS�����_�����4,ͼ�&'5mC��j��I�ג��8k��C
 �4�K�I�+*�Q@b�͑�<�%���0JlS6�/~#�g`׵ ($$Cm�]/������aC�,���\zt�(�>*5�
>��|P�H� }?�A4F�;,S��T�p��շ��r̵����U��ۉ��n��dg?���K��@F<i�'	cdt��q2 ���H8Q�K�lF��~���Z�A�a����[��<���lZ�՟*�;]�;���
���̩��+:��ɮ�)������h�/R�?���po<T6H��܎j+�Sb9D��p�z �r\� <$F.�C90��f��}�A*�G�Y��ܘx�H�V�8%o#u��~I��ΗeiQ$L>˳�L�<����")U�ٹol��D � >�~+�;���2�\ ��܄��7x.3�sF�@�6'����Ջ�'�een���Q�ɩ���Lo�*#���C��a�ÍZ��M�!��+����<��D�֣� Ji���|�x�]г����Ӵ����GF\ٮ��g�7Գ\/������Ѧ�<�ĕ,�T
�7
2�+���j���r�!?����A�a�Ļ��Ff��!]�y[$�_@Uv���󒏄W��dhi-^ B�Е�j�X�����p���˲�ϩV(g�{��r�������ld���p3�l�C��R3�h�&�5���u�L���K��Z�Y�w����k�$D���F:���1R��-W ��tFCC�]�7Q��: [�]��^�])?�߀<6>ؕ4[��R��:`D��� �w��}r��T�g�)�{9�6tB�M�9���b�!Կc��<G����@7��*<��\0��9��u�P�?v)�;p*`M|���+������4P��'�����O��6A�7A����<& ��l /�PSg���:͋q��T"f�dvZ�7�^<�f�B�}��N�h��-���&W@Bn���,?<G�T����f���N�i<ف7��%t�o�n)c��G�aVYW�P#:�j<	]Jy��F�Z=� �M��� ���ݨ1Q�`0�1�i��"\\*ܙIR���M�^�HJI$(B�f¨����"�)�S����E�O� ���8�բ
q��  ��t�ˊ��;b��G f����	���2
�O�`�X�s3тt�r2�.�֢G�ՏZ66@UVMU��%��\-�+���&,��![�b�vll��k�r��25���:{�芥�Bv�y��w ��M�y����^�]���4@}���#/��d vO�Ӑmྲྀ7����nnn���^?�g��d7 �����������7��s1�B}b��Ș���i6LB
j�C�� ��1�f��")�F�9T���1ZG�K�ٝ�b�t��������H}��cz��
{�d��f�{�%Ȇ���,�%����ᅊ>���.��� �ʹ,Ɵ�{��f!9O��]����pD\~1�#�q�hG�� ���>)1X�p� =�C�3����L].2�d�b����{�+�w ��m�"��/3��Q�������p���"�n�{�Q��w�s]�����DK/�Fb��B����)�b�p~�W�ϳ?��=.�����$r)�3p���q0ρ��H�O���.��lDmy���1}�)7B6D�R^�=7�G��s ƫH�&i�&x�0���Jv���y��[���E���2mT�F�i������gpY7���Y�C3=U�3��|3�%&:�v�ڪ'�7�STڑPi��ũ� �d~�-�=��[D/� �n�-���:��ބG!�\~��
���#��w���堁<ؗx�sa �-⓳�&q�X[ԭwI���@Ä���ld1�� !���dr4.�ԏiD[ ��)��g�Si_<=ۈ~��i�Zb�q�Ч��I���B<o��9�4d�Ү<%�M4Oi}���̞L1���ڑ�"���R�K�W�}\�yt����c���'Rw�t��<�Ҷ�M���zr��SSW��@Lj�8Y(֝����)���o�N�>��s��BH=˩-�o�L6$�+w߯�獴��٩�$j�~�!c��2��`���?��V�0�*"�'��� ��<s��U%�2��b�2
�AZ�Ԛ9�]2��eh+Y��f��)P�UZ������HHS��Vcv��8���� Oz�J�)��h�����-=ν�����nB.ń	����\�@=ٯQX����!��eL�iJp��;M�$$$�猛
���d� ��oȭ�^�h9>Wf�ۡl����L5�ݏG�)�25#�q�C�6��+��f#u��-�K?�(i��(���گǹ�Y?7O�q?���~�L�x��aw�	��dc�?@a0��C7VSs�F!�w1�����Zm%IH1k7���k��♏L[�؞\o{�Ԧ�Sџ��(�~���ȟ#:o���Xʭɛ�FO"��ҥK�?�0z��}\Q�����-�U!�����+?O����O�#f�9�Nȩ�"�pYcK�)p��c"��q�G	��tP8+++%w��p���s����@�X[[+5\��z9���*z��P6c�;-OPE���9�N�����d��H����>�����˝\Eu������ +��1�6�멹D7�O�@�BM߻�"�U��}����=g�/�ꛨII��gAg�s�h��ʼ��X�([ *��ny����f�U��Ǽ/�r+���2��_��2{n��!�=!��3�.��31{U�����sz�����'�����2\����$Mv���M��$��-�ꀿ��-�|F���D�)��V��X&��A��?�0K>B+0KrcH�=.����oX�B�ܟf���:�E�����1j��'�<uD:�^���P	�+��.����G�?񳶠R�A�րD
&�6�a�>]���Gd<iry��U2�ʻ��u}A}�fȵV��!׆so�@T|���n|]��)���lFkk�Q�����B��
E�ǫ��w�g������R=ryt�����ޱ� �I��ы�ܧ�C]�0�5n��:�f݊Y���mǾ��}ll4��- ��{9��ѓ��Ӗ�F�u�`���d��1 6d��
� �ۄӼ���g����e7��Rm74�F�.A��&p�U$�9����g-x�(�w&���N�E����`�TG{������x_��"���p0��]���G�r�D�ݵ�p�>y���A�om���s�N�[ԊX'\i�\?rTS�կv�2H@�X��.�f���k�����#�l�3������^
%	���E�����>�D��Sr�F��g��� ,����(��������O�"K�A�ӵ�V@�>Cں���?�-��Q�'!;��@���#��5:hM��	�}��g��,'Jd~��c�������_
tC&�.'�)���	�����e33JJ�G�㍏�_r��;��p�]c�?e{m3 JS �p����D���J� a��@�_3F֢��6v�6��������Ϝ >%桫�U�xKe�#G�V;ٯ�b�I<k�D7}qz��q��sj%���������X�+W�dH޻��Μ{� hɍ^��0�R�1[U�ͧ��q�P���'���b`��3>g͂�z�oɓx{�E}}�Ҁ�;}�[�.j9��}�km����w�f���&6�����V's�G]�xP��D���<\��o;U��]��!9����Lv��v����[e�+�o4���}�!�S�\��lE����g(�d
6%�?~,��+C)���'��-��󵩮��]Ko3�A���S��DT��Q������bѦ�"2�	wO��ē��a,���3a�#f�)J9���&�����A�f��΅�ׯ_�?'X"�bxB�K���y�Z�7PnK��5����+s1Y��X]���{)`�<^'0�qp/��_0r����=�(�V���ݟ�i��q=���7(I��c����pw-ޠ3�k�v����>~� s�d�BNT�K���4�{=#�3E���TWdP�)^�w��w[�C��K��X���I|�;�Aҭ@O�X~��vݿ��r���s�6bR�]�a��F���:�#&X�'����qG�RXҬ#Rr1��Q���(he�));i�5��q�kޖ�R���h����[A�]���� ~jqڸ���Z|5#�[?T�HO3w*�l�V��6By���3�)o:[BW�om俼ə�܄�	�U&�j%J��.�bTg��un���R2�=��۷oY���l:��[R�Eﮍ=�ä�u���96!�}��(��}q^����{�k�{ON��b,�&-wl���7���e����{���y��D*��x����M���V�լ�F�5H�Q(�����"�V�����T3�"[!)W�ZZ���K�G�D���@��~�B�n��T6��CRR���p�ѡ(����(|���/pa^��0e���mxEo4�H��j������Y���+g�ҼId������Q�����,��W���9S�,��-��g�3�T��J�)��*]}����!Apq�s����Ϳ�c���Z�|)�|i�(����&:�s�,��²�7J=��eW���ݎ����}��߱W�6�����A �&h�6����X�!*<l��.�'�S>���rc��܏�lB��IO�=����D����a<�z@������ӑ��&�H+@�ThӇ���[&�RD�8J}$YG�<Оy~������=��J��/��qy�q���J���6]}#�u1�|�$�T���	5�'&ބ�`<ˊ��Mx���ڜ�G�!�T	,�����O$���7�1hΐ�_��T��*=a9���+x�� �2vȈ~����Z�Rut�8��B���E������'��}lP�N懺S��G�؎pL�;�u�Ol|�����A��7���v	hh��(]��c`�	6$����9���%NjrU7���B^��7OU~��qN�'hOftƀ�̪>����]h�N�;�6���F<�e�rf��*���0ʌfh)�w�R\�¢RH�$�q.�Qʸ!-'�|z{(��3���6A���F��'��Oz���z)5���K � '�YJ-��;8\U$`�?��Ml����ZR�K�<}D MN�i(lxX�`S�y��`�`̀���Qu;�f�i<��Z�H������~7"<|r���]�3�E#�}TK�`��[��⁷pt��4�b��i�H��.q�����(Qڥ�0 ��r��1��C�����:Gf�'������S����R��O13e�/Hf�����+��/u�G�%8��xυ27f�@�tmrU�7{Xh!��0�,T������<��Vǅ�����Ȏ\(�zC���`e�y�O|���V�矶)ڲ3ߵ�k�Kwؾ`T�/�#��H��}�3����� �F�0x�>�:Ǚ�u}x�G-nM�Y�8G���c���|@�D#�In�/�zT/�*�R�DW��:'�_9�fڗ"d{?�n�S��tݟ�-=�R��������J����(T�aL�q<��r�� ��`*.�b��(F�-Ne�������Z�~������)���T���_&��i]�ϔ]��t� ���]�(
�����Ng�S��<f�Ԗˉ��o�̊�<�����T���rd������>���|��4ہ)l,�1T:��P2d�Lp�}8̧���'�)��Dm����`a�m�s=?N`;��V?��tCSE`=��K��2��Z�-\/�`�GZZX��U�{��%4���Mx75���G���eB��_���a�Ӎ"*ė�,�MR9�{�=�ɇ�_�f�����=��� ��p�?�s䨇}���׬�\��Q]Bm���A���J�W�c	�(��p��wa�Ú�8�-�L�bצC��W�\^�
ag�ߋ]���ͽ�D\�[��{���#���o�ǩC����7�8�tN��k*k/ m�d�H��dPs�*mH�B�H�6�χ�߯�uK�=��Xiz[��c-�6-���o�O���n�G�E����Pl���؅ �f���c��<|/��Ҥ�=��&;��͆����yl<j�뽵�������۵3���{B�03#���3��h�rhĵ=HA��f��)n�޻���b�uo2._���n>�_�5H�QW��C4v՚�8U�wQ/�9EΫA�_2Gsd��~l�_a V}%���8���#w����@t3�^��7�]%�5;�H^�b��3����'�y`~>s�l��FF���#�HǑ'F���p;��5c��o*�1Psˊ|� ͅ� �+c��'�@EtØ%�n��Y_�ڭ�Eaa�R!]��Y72�/ad��aέֺI��1��T�����o��^�i���x�%BY�s4��b�*�q�*$��A����jQ�|�;����'�0V~�!:��s�����)4Y��հ�6�Kgv5��_����c2N�WW�c���S7�d���}񹔆��\M��*�I�Zq�w8%�=&iߧ�?�&�w`��R�e���XA�|Sx������|�]c]o|��/�.��ϜP��ߢП�gԌ��~�m�=��߶�R��]���ӟ���"��x�:��|<����'iy�(48������]��������7��&����
�AbUX1��Y`�=���!�^3�v]�SB�?bD(�&a(�uf!���Vc�+j��a3�H5���U	P��l�p��7�'���|VXHڃc._ׄT��_;y��	��[�%�c-
�}Hۈ	�/HwN%d%�N���0�q�`�y��NK%�e��v����N���<{�����#2q�?�-Fsb@U��(�#�@����}���l����ۜ�n�O�	x*���%yfk�֬�Z���Ϩ�� �*78�Îb�<Z��i_Ȩ��h������k���8�Fq��3`��=Y���p�����R0��갚�ḃy
�ˌ�]W�UT��'!�F$�.��.�!D��U�9.��R�@ڗ����|��
�|����Ӽ��_�>��{_6�nk���j���	�����:A�1���N��_ nK��=����9y����F`;�^`��Ⴔ�B���L�o���՗�4�$�O�s@q�뒵���ꍂZ�%±�0���K) t��WY���R�F��'����������,�t�f�gL��}ڬ��6�6�Є�)��E��
��U�6�8WE�}���au�����y��fMě�l4����/ƙ���QZ??QD��, 
���]���{�L�q�����>?���4v9X�ɝ9������SK��+n�x�a
�d�嫯)�`�r��4�2����˶�ҙ�@R�J����:���������~Bk��(��<��洮����ɯq7�%�vR	�3K4E�c��N��؃�<�U�!�=��M�/���U>9��w���:�|_瑟Y�J�y��l��pw�x���ȓw�M��&�q�~�k�B�����Z�^�m�T�3K�*2H���Z��N�9��u�;a0YN���8���s�s��¢n��J�ez4>}�q��ٿ9*N�xP���*��s�{wAe�byܾt��w��r�bk;m�G����wZ����/���Ο��R�_8x�V��V�q��Z|�N�K���=U�����/�S�oWEF�'"�X������̞Lw��|*ӥ)u�/2+Fq�ǫ!��}�ǽ�z�]�c��AU˺qK����ɒ��3ݱ��нR�u�}�π�7/���]���d�mՁq�c��-��=k��J�٫�5h� ���Y��r$TM+헿ךlƨ��=:����=U�"�n��Pem�p�
1B~�x#��Ke29齙�'��~�H,�V�Ԉ�m�D�	��e�_���Q��5��)�%���;�0�� (��d+����줯�K4E�0��S)�Ǜ���Sw��h����PoI�v��2��#{oI�ԫ���*�;����mh,'�;�S�n�F���lM����՝�ӖC�pVpPj}/Ų���$|a��(}C/'B�؈��OH�jﺾJ������G=0�3��Q��$�zz�]��,nN���R��f�Og������DLC�a��A�ԓ��̡�aȡ��&]����C�� R�����}^��#�����Vg��~Tw��W__K�V�`'�?�>�*r�%���n�M<���p[$��w2?`�7E�zb��`�|�������5P�	��l���bu׷A9���/�$�?cʡ�u�^(~%m-o��6��������%Ѫ�8F$p��*$�|18)h�_�g�Jav��C�Vi~J.vR��7f*_�G�su��ڻ`����s��/��
�|1���*���Q���@�k�T؍��TW�p�W��g����?mP>�`z�y�Gڐ@B�_巣`4���Qۃ�Z�;�-:�1/z1��p�S����JPK%�$�!�������������>���M�W �F߸�����ӡYS���%���":7]�~���>�f찥��3D,����ٰ,p�,@s��`��_/�Vc��%����U��a���Bs��Էa�r�d�c��絭�#�F��L�ۧ��G�2F���
-� u�}a��<�P|g,|AH�!�Ɣij���6��ĉ��V$��]��<6�.7 *��N>��k[�c5,"�u�n`��<5�!5�o�����<d���z�R����P|��8�Ɲ�0���N��$��Q>��z�&.�o/߈�Rئ�'�d,�u�>H+���бƮ$�����^>cC�m̔k��p������U-�,x�L��b��q���o�A?g�������юh���,=3�'`��<��O�ϝ+E��J�,�+[{|�������V��xNF����Gm@����`u�X��o�)�m�����&�P_�,���`�9/C�=�g|ݸN^C�������*�-9.,9$��,������W��OE0Vc��n��k��4 �ԓ/��	&��X,�W�*�r���뻗8�oYG랉A��UBB��V-�#����˜��S_Ɠ��oS�)AH'���Ig�b���O�������`�l���;r�7Ի�:����m�m�:V�jQ@"�ٌ���j��UJ?>n<\Q�wy�X9�|�&��)4�!��2!mw����fO�G��}�����UC��Coķh��Q�mhj���[��s��)`��N�tӗż� �s��OFE�9p�:(�������l_{=�F�?{���_�<�s=s����j��&���R,�#��s��6�ثAM�FEk���"(��*p�p�1��~0�7+d\a���u���������p���*kڂ(5��m��J�3�#"~��?~o�k���ŹXP�Kŀ�Vc���V�fm@���'���Մ�u�@LK��R>�XԻ<*�$Zm��pX�5T��ߢ'm��y��w�B�1�k��²��⓲�ǯE$DN�f���7K
˸���{[/���6�ɝ�����om5��6tⵌ�Dm��*'�K�ޮ���jA�0�P�Ju7�,��;Nq����P�a7,��ȖA�Oٻ�啘�i�32.�����;z��E1U���]X	��������0~7u��N��2�*��{���A1�?o7d���z������v�/�;�h+���-DՌ�"�ޡ�\IG�Ϙ�)�O�j�U7<�j��@K�R!������T'�R�-�������X%�D��][�����ӭX�T4��Y�/�M误u䏓Q�>o^�U��X��vS��h��~���I�`Rt�w�g�͈���Y�����/#�3ƿ��wMx�1Z�����nCF�U�9p	k�=���Zc�Qܺ���ZtR��v�:}Cl��d��4��^_]�Ή����D��2��?s*���֭�Q��9{;l(R��Y�����#L~��P�\��1���%}���c��+�c;:	����/�vm�<d|vC�(O�8�t��˪�&���!���(��B���>�"���;$8흩X��Ŕh�缉޳�C�;�Y�g�p�D���G��V�������O�uy嘘�:,i�׼�䓊�bAz��6�ڿ;84����6�=�*��D>~�c��d&��p�.��P��a���r�U�!~�eͫOi���5Kb������CY0P+�[I��B������_=�U���*i��o�|�pV$���º�L�b5)�Z8Q�4�Vu�z�f�8]u�*�q\JP��J�*�}�0�\K�O0�~��P�����O �qY����o�W+��i_�ܜ���:{ ��mүуL�P�Tx�>�]�0�s�Uf�P9��;�����=��SS�|����r�Λ_�&����&�۞�]�]�l���,�z��C��ɒ��� �͐g��C[_����X��{�J���k��rwN�&�6ė	*��n��A"J�Z#��os7���jy���\�t�:�c��_d���U�-���Qo��fjLP����U�XA4+[�q�Y��b~�����qa��'2h�Ġ�ܻg�e���lY=EA�2����F-{�lZ��l���������w�_R�1�3��>%!�6SE�"��ƹ1���ua�>�xːü�_�3�-;��s%4w͑��1������P�n�}�CJ#~�1���R�E�;�>5Ξ�n}��q��"eK˄�eF�͛�Q~���bU�^���/�:ho�u�p|�w��zk�E���q�a'qO���ɬIcnQ?����"��q]3��R�)l�U�׈%�hD�����V��L�z5�ŧ� ����WC�pZN�gN�М�g���R��ɭ(Y��ΗP�_Z\%.�|"ehV�ST�t8׭��5���~��\��GI�����:�_���Lk'�-�LP>z\ɖ�9ob�D`��/ף2�T��9�:�h�=��ـp���e�z�n������h�T�G��T6�q�̞HY@���jo\���}�����Cv��d�x�.�d%1��S/OK54�$�����G��3�\����.x��y��ͽA�Y��w ��ֲ��US.�D��s�f�?���X�;=����o�0��	��׈&��F�����N�T����@�2�NRt����͡����/)��9s�
��&��Q�u�ǽ��(��l�8��t|��k7��������]��_���ؚɂ%�b/�z?�x���5�'9ƞ��w�N��6n֬;�FZ�Dd��\,�)���ʠeP�O�����^%��SCbڜZ�`m~���r\Q�(.��l`�b�91�8���P<$%q*fz����G���>��QB�*D^q,�M��<�$~���ɇ��R�D&��t_�ת l�2�����mQT)ۅ�u�K�e`AUtQ��б�χ�M���wR<}������u�tZ�[+��
��s�JJ��D"�r�?�0s��{�>^�/���|���,^��(�{y�?���F�H�M������I!���������\�i�h����*��;����N���(Rk�'��a��_��0ń�Ft��t|�8��gz�V)����(�aa^3��mt�L�����]��B��U?1�-���#��%�PoY}�{��6�cOQ�/�41�f�Ǧ�ecg��l�>2j�Z;i?��WqǓx���'ٵL<� �U�e+�1J�K�T���R�;D�Ƞ)-��wF�Z+U\,eMd֏4�_8MV�)o��o�m��� |��!2��ߒ)C;eP�®�k�[m,�T�)3�V�6�?>�y6�3vA���;���܅�ѥ��*�8�^�5V���{�;��K�	zП�n��u��y025���/V6HvƿQYu�����C弟�`N����1K������,I<9���|�z�����w�a�(1�ŭ���vy�d����]o�'R�`�k]X%V��%�JQgn	�#��U����N�l�����ܢ�ء�<�JfE����,��L��"�h�EW��@���9�pNe�.Z�j65�ٖ����:�I�R�����b�ȱ�����[���O�ڤ��y�L���E�~���,�h�N�N���PR�{��Ĉ�`������Y���7��qUV��{w
b~jr�
���u��-�i�:�9d�.)��+����eۈNt���Vqvtnw��V�3F�u�=m`N���Z#��|�7\�[��`�X>͇yWMl��0V�9l����t�M�g�r��ʨ��O���0'�)W�j��v��\��M���V�/�(��<ȃ$M�Мq�ʥr�%�U'�s@�%��ѣ݀�elˏn��,9.V7�z�S~L*��O�_ �N׌vo^+5Aw1�k���#yS���wh6���	�9_�ԕ\�u�$��o 7��I5���GQ����+ 9�QrO��ڟ	hH�}��/��\��x��2o�� ��i	��j?d�u���X��%!ɚ��c�p���>s���En�0��$8N�=�M��k�[��T��>�쥈��×
��m]�)~�H��ȑ�~�b1O��:˱�����>X��8����������lf ���{ϰ(� \E�EPTT�
"�!LdQ���$�!��dA@�"   9*I�HF���3[���{���{w/�9g`���ꪷު���\&�ڦ��������~��˹��
�'���W8�O�RE�ei�tI�ı��]��g��ʝ��^e�g)ݫr��+��gq�d��%@�C-����5���n:�|�+W�MC�BSV~hI��+6B��@���%���A��Ky�'�+||��~ϟ�^�ksJd�d{z�D%z{�'O����[�-y/L'Vx��2�P�-�y�}��,Ǵߵ���6�4H5Tb���L�$ne���b�Z$�{3R+I!�z�����'�m��UV������ Ý���u��S3�nʞܬGq��Z5�M܏U�5����%��W|�`�v��<n�����薈k���}_��W�3S��<P6����d�VVi� ���m��.��=����h,�����S��W�B�OP;�`lmCU����뫻W�i���lJM�5�уC�ɿ5�y��gR3|�����+�f�����3\[�?ݳ�=r�}���������']/)���[�fh���Ҩ�M���SO���[��h�W��� ���a%٥lǕKvo�V�P}|������k��n<2�U��S?W��s�����V����'Nd�o> ��(��[g��K�9�L_�2���-H$���S�e��i�J�9nm��F���<��%�W^��\���\z֢z��}�=�IA�{雗��!��
�6����Q�z(7��5Z2\�bR���M����w���X��	�Hާr>��+c�ƭ��L >t��FM�`�E��^�k���_G���J��zs�rd �7��-�Z�Oj�4[�<�yJ�����V�Xu�n��m��ʢ��ql�-"����FW����7�טZ�,�5�,�FƖ���g(��nm�z��=9*}C��<��'�i��mO���di�Bj�q,%т9o	��v��_}�"�JhD}`�_��t0�|S�"[��&� �>�+��W�S歼�C�s��2ç=���q��h�+;!�m�����r�����I6�����X��Ӣ�OE���|`����͂ڝ�RKL3$���O�
��Szn�ޓ!�ם"��[�[S~O��%H�ɋc��'�N
_�M��Y�t�|U~N�]�߉j��;3Gy�;�Rۑ�� [�K�7�6�A�%eu?���h	���^n�:'�5���#�3��+j�4x�F���GG ń��+�5�O8.���������k�o��D2�{�E|g���{wi���,4~����y ��� ��:��/χ L7\�7����J���3|K�D�5ǹ�Ж�gT|�z���x��hZy^�0�Ǚ�u�=��o��~�n@p�͎fhd�j�56�h}�r(���7��}�fRʂ�Ck��e~o�++,}o���vxqP;��U�����ǹgߙ�O,׷����������N�;V%:n����8�asنr׾0���ë�[vd8�����.vd��u�E�K���1y��RH��.�ĩ���*��7<si������wr�I0��ZQ�ڼ���Ϲq���� ��[�4:�}N�[/z/��s�Ӊ�It�dN�*�n/�̻0�f�{O�]ɍ�����
��D��-[6f�F��2��?�>V��'��NX��$�(s�ߥLz�=l�<�6f��#~׾/����zG<|4b�\=�E
]��Ќ���<|�b����Sz������a�ƽ��_9�}����bQ�ѦS7�͟�S�h�;e7I��v��;�O���^J����o�K���͙'�]X��+���?���S.�����H�:�w%��;4J8Q�?y�|���ע�!�&X�Lh�o[!?P�lq�C�Oݏӹ�'�D�}J�9=��</}e���w���}O�};rY�e]�3��l0��Q����}�ޘךϔ�KZkr���Nq2�_z�p,�߲���,�������	'�H��>�]s}��9��[����W��W��On��sU�n&m�������:�g�K.�,VtF{�*01�-Ŝ^C�Z�ރ��5�oH���O�V��t�|�ؒ�woU�>�c��?]J&�=��d��|q�pCV��v������_�z�L�U����l7��&�]�!%ٝ~_�������+�ϾԴ[5�mE5`���뗛��ľo?�m��Ή�į�*?����۱:xF�髯��"����Jc�e���ON�#�������}ږMۙ<n�\:yl#��MΒ�y�?]�,f�1��ʱ͗_��sYS��_1��s�(�۶���fP�N~�4L5��V]�RH,�7,<�����F�&���I��w���AJ�geVӺ:�퇍i½F
�%
Dw$�7��(��c�"M�;�%
��sVT�Z,pqCyKsó�;�N�J�Q�
��J&1�<m�*QN����#�t�~Z������[ڛl��Ժ�R��9���3�c�����LVsg���5�=V���:h|"��zL<I�?X7H�~JpLs�̴\hg>4d�h��3Y����K	��{(a�E���M�6�#��b��	�ܶ��_�����J��H�*�����[2�.�ʝZ�d\�M��,�pƑr,����ˮ�+#�������{��������]|���A@E�5�F�hOE�81qo�b,�.>�k4�G9f��{�ݗC�
��R�:��D��S�i�GJ�56m9�1E�x�tT������7SRJ�x9��hIF����S'f����9T����b|�j�S������ܙ�./�/���O�s?8á��c�N��n͍r?����~����S"@a��]���ゃ��*�^`6���
�S�5\���F�sg�<�l�ݶ�j��
5)s�ۖ�z>��d��n�8��c��@���޸����.�d�"��9�C9��?��fi����J�Y8�{�&�J����9	�iŜ���#�&�<-�8���^����,��Plq�>�lyZ�~�H��Z�-�cm�6+�3�q�z1er��Q�Q�������D���T��kdJ�vf�>X��<�T/T)6\ju	��d*&���L9�;�30��ޮf�MC���mU]Z�!�J��}�-������Z��à�Z'�A�e��n�!1N�)�������� /L�9{�!!�^��3l�Y���.'ǩji��2�ތ��v����X�<�9�:��n����Ie7)�����Ws6H(�f����MY�Vs�¸���a�3�}�G���˴^�t�՚�/w����۟�2�,�qϲޜ�&�����|E��vYtC�n˔�)A��M-�-�5����H���]��`�i)~Gmqt7���;��2y��Ȼ�ߕe�Q�dO�u�p�гTt7����	�B�吗�����К������6*4&
W0u̴j��|籤��(I*u���>Q���+vw�^�u�mlc6�� �M�F)�������em݆��w�#��i�M�F��H��U����e�����FB~	^�����NL���j-�`Z����c���c&���6$��3L�LԪ���h/;LFv��z�}9}���g����$z7�*�פ���
�+��O������7�?�4r@�5e��m��N˦a2���]�?M���1�'�u@J���8Q#x�;[�}~�5�V뇅���WW��R����$u�:yTװ°yOot��^��-hL�<�n��M�Gh*��d��-n�[�Qy�o����>
�b0�ْ+4�B���@q.p�e�g�=����[�lI:����c��;9�i�bI�N;�l���������P�tQ4҃i��$oF��_'��~�uS�}���`&���Mf(��{;���P���gϲ߾��}�t��g�6?\X�L%=%Vkx�e��Ȝb2��r$W�s�G?H�ّ�2��W��'M��i`y����!�o?��3"��?������$��Ӣ"�5�R��]Ф��]-�nl�J=�k��̍�M��d3�:[�4�<�����Б$�7_���������<cf��V܆��P��3���C7Zw5��j�(`�f�d#�N�0{�Շ��֎�*��\��%�J�zu�GD�TFp2�Ns�VG\ԃ��־�c,e�������^�`������6�Qy��u	�_��Qޫ ����{��y�"y��*S�p	Ec��g����7������(�?!�yg�-�����ݯ�����+ct3[H-�Nw�>����^Pʗ��H\"MńgK3zn#<g��$�#��ډ�훇�=��2�6�����!\o��f����*+�����;]/^p�1L���53:���4Ϛ�:MZX�$�D�����	�C5�	�Ő�6�)I�_�A�~��&�~������;Z������I�؃j,#�:D����saN�V:9����ī��J��_�d�|Wj�2�>��mԈ�E]�~5�g��J�ͭ� E���j�ڷ��Bݐ�V�@�|�u�P�nv�k4�:H�)U��G�)�vɐ}��L�M��k�!)8�����st�;Ty����=)�3� �Q/�'V��^���gk��q�B�L����P������|�iG6l��oQZ&�~a����{����w��3Z��;��fw*�i�Kp�Շ�˯��ߋEI_����M��F-�]�v�)�mF*�Z���.�0�T����g��E;�?j���|cMgǴ�ˡ_�5��>E������o��Ye�33�H??���l�i��5�xp �)����?_�F��g*�g��rMp�;�Ln�d�2�MQ��z�&��|��Z8��ģ��ޟ���	;�w����ۆ|`�ܞ�J�d����E�]�_��N��o�������]^�.�O��'h�z��X��u��"�E��\�.r]��U�+Uq���|�xjP�g��G�{~�����O��?�Z���i�����O��?�Z���i�����_rjLL���Y8�q�s{���[g�Pܣ,xGⱑ��wS��iՅ�މ��ֺqqI&{k*=��:��w��S��������T����x�ߒ��~����,��������u����\�.p]��u������U�G�	�#�b��ȓ>~��ӄ�F���1S6	�o�"�����y�>��t?��(&�md��]����2�8,���L4,Mx��Г�ݽ83S��}Bȫ��S�P�|7�͓��V�D�i�H�Ȭ�Z�xTEO��e��,6MU6J����2U�`J��l��ϯ�eU�.p]��,0�?��]6��5��3��RV�%�Wv�;,�\�������̛%�/�g�_�5�1]֤>�g��1�ǉy�B�sU��|��ݨ��v�8���#}�������Y�����br����ݪ|�̌q��k\�.r]��u��"�E��\�.r]��u��"������ �o��gb���Lmm����Jm]�%{������a[��Xm}}����B�b��*�鮮����\	�� .��� .JJ���>~�~�7B�g���.Z�k^����7 i�E�8w�N�g��[{<<<�~~�/�����+./_3�0??��cPa���Ϙ�(� TTT���虐�p��A75����t0��9�����c�߬�����ի��������ׯ���	��(��������S��TWW��:p��0Hx1x0Ix|~��k�g��h��ٟ�;��6 ����64�c�>��~JN�dkk�)�>~M}�%�RU�16߫�||fff�x|���,�4)O/hβ�A�@����`{��A�F�mҮ`�dɻ���X��U����xCMMm�×l��zz.h13m�LG;[��LgG6fZ����[�.�|����Naئ.�677���:WVV����4J;r��\uһ�����V77�y	�_s��(l˶�
4�qiʹ,N�(ަJz������6G+�%�oJDC��i�_�	���6h�52���mc�\�|�zC�J���0�Iǹ78˸^�ձ�E�8�=�N�Ŵ�P�z�ko_�K�Y�~a=q߫����9Ϝ�S���f$l�^$��*���F2���;������LNM]266V6-�wI��XwE ���Ru{;�NU���쯗ҝ1�9��˳�֤�������bѠ��jN��ąߎ�/�"*{3<3���ٕ���Ƒ3{Tda0�1�XVJ-LzI��A��(4K�o%iK~������c��Yk�E�Qk2Zi�%n�p����%i��;���'t�PʹZ�M��W�+Oҳ{�f�:]�;Ǌ�T2�[���������E�|we7ڣ3]����08����}�+�|�����HfOz��8�aw/�ypL�I���;���8�v��0r�`�綱�Wf�~v�|(������ܯ�cs=���C?��O��_}xT{X/V.J,Vh�Q���Mu�~�Myy*��8p�?5�;�F#�+9�����9b0V#����{R���J��A�R����;ev	d�SS����`w�s�����
ܙ�ƽ�lmm����000�6��Ps�I�#��->w9��ʪ�3���B�.IKKM��'��}�9���Z���M���y(�Z�uHPa�����M��1�XĦ}�&�)5�F��^�����lPs�<����N�3u���D�#�@�g�/^����l�cӕ���_/���r���$�R�ӥ��m��$iW�N4���S�u�x��2�\!

���ݢ�q$u�)_��:|����:Щ��S��[�8Um��hU��
�ۼ{�K��D�U�@��/O����XJ-��9x������0�Ϋ���p�̞is�M�/�Y}z�����@~~�i�$�>aR�y�����:E�C�<�B+����-a=y�5�>� >���f̥*x�aa/B�ͷ���vGQ�F� r�h����;�[Y�e�������9@R��?������W�up�r��������E���B�-����Ѐ��{��"�6�܌A��3��%�%��m�l��K�Sc݁�E<����09M�c�8�T'I��{�޹P����~j�����n�t��]O�I)��;�S��F�!ŹRX5���l��v�v{�j���6��h> ����۪h��w���?^WSCe�=u��0��mߩ�.��.Dʫy')+/3������a�f�,((�D��(L/W�cojty�]����׵�/f���$�L��E�~��m׽`Gr��gQ�܌e�ٶ薍ۙ�xf"�>�bͅ2��M�g�n*�,��aQ�U�/�� ��5ި�}/��\/��լ)�<��}%ZN�%JS���{�^-YY��'{����yfݞU"FE=�^%Peq�����~lz}f�UKz��U�I�<bo�J*I֔���i2�S���/w�ªu@Տ���^�����ʤ4���["(��d���0ĩ_�~���ɉ�*�;��<����[�@���U��l7;
_��C��i7d��v�1�֚�TΠM�)T�!�S[�o����H�L�n��lsC����vUH�fnN�Ѓ�O��M�T�����Ӹ�t_��J�����/؛��h��S��~�	KN��ne~��}�>U}�1��u��ϋ�/���ܯ�<�����:��-���E�~��=�2zʗ�Ҟ@���:��J&q͵��܁L%��k������A���wg��g�s��ͮ�Io��.�ğ�*��2�4����e#s���}r����eذ����.�P����GJ�7��I�
�lŷ�$��N�|H�d��@��[�K�DO
���:��{�awF��fy�WY�#2��^�mMK�b�>=h䬔���s.J���fө:E���Ϣ�T}1�3�m���O[��
��i�%�?��D����A)��1��]<��ͷr.������k
�݇��-���ݰY��~]<��(�L����8����Л�n=�[2 �w��st��9JcnaQ1�q��݁)� 0S	SR&X��!6&&�H�k�>}�$����tT�[�y������8�{�bǁ��+��x�F;f��r�U,nd�~��D�N����%D�_�CM�rvn̰0@�l�˫�JZ��Jh����� ��>UZ\jJJѷЋ��e9�Z���g�W�e��/]sS;��h�X!���������xR�COy�PP��|C�H��t�����奅�.���0؍~nL3�+�B����Tc������T ������_s���|M-���2u��v�3�ť�{����_׼�	s-+%v�/��+Y<h��8�c���pQ[�WL0�*�R<_{���tg½���+���v{qU�3U�F��gZ�4`B.O*F��8� S��������������0����{m��������� �3#UR���B��Ϯ| R��A� LT��J	�Ef���^�S�7i!R��2�a֨�▆{�5�ű[i&������3t+o�A%�7gy*��������N#>x��T����S ��Jݠl&ini�g�m�.Q�E�mA���75�:tȴ�`Y�'��;""�F-V�GV�ԁS�kW�������$��eO7ϖ*�xH!)�5�NO	��Τ���(A���3��n4�K3:=��[v@�ޔ���˪}���v5�bl�
�H`�≛q��v-Do���]�[��Ew�!�
r�����ٹ*G��ed]������N���u��ҿ�{�8�HU!$4~����X����%����o������
^�n2����:ؒΕ3�a\PH�F�,+x%.��N!~���*q�hk��X�,���9�KDx�xx�bX�g{�)���O����R@zh7b��v�#�Bc0"�x�|H`��m��I)m�:�A�e��:,��?M���N�x�������w�oލ�9����Y�,�3�M$��Un}x�G_��hG���EE��*-�u�}hT������b@�^J������q.��/Q�8��)���W{�oOň�瑟�A��񘋴X��}�<]Qg�[ס+	l���=>��ZG,���5#��k�E���<-5I��w�\��;s��M�ԇ��vghR⒳��Ei!5*�d}K�YE�.��*v6�WT����wZ�8M��vק��������J�����d����-�=q���~)k�~�m�ɛ���� X�|mꢽV!{��JA�7s�� c����e��vl= ɢ9~��]�N���(m�;�l��2�@>R�#5{Ȱ�vu�QZ@�sWv�%c�|��𸡶lfٖ9��u�MY�Bf+:_���z2ι���.2NŬ��Ӽ�� �M��I(
�D��.Ͽ��tu��Mo�l`�\�d��m�:�%=N�g�}u��+�\*�.�HIkf��Tٌ��7���yN�bQV����1���-������b�W��TLuM�K��_��;�+/�V����VU���J9I\���`fG��ҫ��4�fm��0<R�h��0�N\�BL�lc�H��(T{�]�i[񯒗0�w����|����"M�h��-�&ʹ�X-t:\�J$m��7��!t*C&;�w�}Vܮ�^R��O38��P���D5�'c �A��#������h-�ތ)�]��[xȲ��Gc�����%��<rC"�������ۗc�o��pRU��$�~yJm�'geiD'�~��P���!�6qo�򸼔���egl!�F� ��WIJ���Lt��b3�*����0��r|�u��`f ��`�9 *��w��)��4�R�� '�;
;��Y�"ӻ��R�"WE��g�۲��"`���T,[����K�<���Q��^��y���N���P�R@����=��J;��`�s��~a����{��Q�f��kF�����6\:��[�Nh��>9�����s��JP%��������^�u��寉!22�t���B�Q�M<	U-@<�
���|�e�㭳c]]����$y;&^���ug��� �q���s�A^M��V:ƹ��t������kz�y�v�;�9�^�u~��{,8����B���޾��+<���4@�$��`��.>��� ��Dۇ�� ��J5�~�WV^���*:?����]�\0�{i3؎*�M�Q�ɞ���f�7���X���o�%q�y0vW�SE�NI�>�cjEح\{<��00~�#�E�4�W��N!'[���Z�N$uQe������
�Ri7��^Q���/*�N@�8����Rǵ+��I�B��1��Z����dM�����J��������:��eI��d���,���{R��T��a�1*�%r��3��8z���/h��g���l�%�m��ݹQ��q�0�1�bL]�@#W�L�Vd�i�j��i����P&j��	��({���B!�Xz�=�~�m�U� .�"H��P������`,,1U4'h�}�D���v$�02XS'R��a�\����91'Ǘ͊;"{K��f�H�@u��2wA/�;��z�6	�d���혧`�{]c���I&?��J5ė�E��I>��.���r����΍ahq����Cy�E'̱�xGP̉����>i����!cG[��Uq!rB!0��*戹�*���Ҳʐ�V��رr�*Mj#�I���W1��:�iy�`Rl�UK�by��֐I��fMF�I�r���7�m�թ���Ԣ@�:Ss����:��%��?Q��jɣC6�,�b��)�b��<d6Q�WiA׶�W��[��"c���Rx�Ĺ�?�{R欗��-;�WU�,-���W����@{��t"f�V�7]��Ѿn����2依=��ږ�� w��pKz�VV�M n~�������>V�6[ħͼ*��/lYo�ԡ30�Ŏ-M[}Z�!�'rm���)z/�f�������TȀ ;t͏<����`7,
��e�ܹmܜ�1߭�����<�2x�|;���~U���V,�j�P�����3�$ˤX�c��!4ю�jev��*�����4.��� :u}��*���;.̂�6䦂��/ʞ�6H���>�|皟
$Ȧ/�bn�:ʜ��:��L��2��k�Ɛ`�~�'���O �*{���|+�����h~�Z~���A¸��!�^x�N�}�, pX3�?1�>ɀ|�t/`�vz��s����W���	d��@�"ޡ�]�UYH���[OHR��I��⡂8��THJ���!R �{�.PE����hs�%�t�K�X�y��!�VP�ؗ� U.q��Vu۩�=�
ZP��)~��%�kc5��ܸ�3\��X��G����s8�}�w���Pk&_�%�E�~I���NNN�T���Sa�FaV�)��>�Kj�@���:����H����8A�8��_%0�������˶ ���R���\��?��S����}2igU��	��?��K�uvX�/�y�'j�Ĩ�|��H�;K���+��҈�A�����&���VL��Q|��ҡ���]��o�b�,D:�j���`�T�?���W��rQ����d����mY�_�ì6�S���)���0�0SW��뫫_�ri��5�|�i};r�z*QIO�������v�+֬J���Pq�|U6pv����[�+Y
�0�����P�g"~�#�v�0Þ�fX4m5iO1�`^��[���n�Xd�)�x=#����L���_/��*@`��ǻa�Ϊ���ޞ�a^�:
�f�3��[$l����\�Ji^��,]���dMt��{�˫J��g`��%:�����:��8�@�gF]7"��c��xh�n"W��� ��}�G��^ù+˫��"�Y��p	�J��9�^ ��y������}��$o�
A�3�QYe��A𓸴NW��_u�d�`'_�s����� �
=��ӟ@\������9J�/�*�D�sdϴ�9�P1=?r1�k�rAA�D��׃E����ag(r�#����!�Xܥ�Оc�ը��_�iE�9�ҢJxF��:�vlQ_dp��l�C[�T,)$���F�,����[	GsH>�/�T�R2��%���a�79��A���.&�d\��ᩞ��=O�I��:qC�_!2�F��(�I2�qV�q��zZ������ TW)�e3-G<1+�V�d�ikֿ�n4:�fړ#�8���0Hp2��O����P��6��|.�}�ɜ�zs ��+�#+�#��rK�P(#�c5���%Q}G��F��Rs1���3�h�JZ��,;��̫W����Yє�M{�D�u��ϪE>��\�3]+�щP��+�'Nlt˟q䥅}a�Μ�a7T�]�GJUHuG�X ��Mz�Z�&Z��E��`��m�#���섩�I�K�*�Q􍓮K3��S��o��*�ܤ����I�Q�$X8��uG�y�w,���ϴPi���rR5[Y�Ꜭ���x�TwTd���A> �|ƪ���Ӯ�B�w���?b�d�;P��;Z��
˃�zy�*�X
��]�����`V	���,��皶�9.�a<nu^���}� �� 6Ѝj�qqq�;zy�vxAz"�e<�N#{���2
�H�����Ӱ��P	j�+�<CګM���T(`p	����n_ �a)��|"��VT�ƒ?�\��x��B����� ��Taʫ<dV�	q�f�/2�*�!V%�e��d}�Y/��� *��ɒJ��3�ˋ0#~й}��o5��]à_P�3Bx��1��j�]��=K+;�����X@"��!�J�	���k9��,t��`F�g���W��SIh��m �92�"���������Ǖ%��R��'+U	��m[`}H�*p[Ѣ�*�S�����T�JƄ�A�GT���G�"��^��}��M��]}�y`���@=�Ѕ#��G��"5�ei@�a�A���d�o�BbP�Y����,�	\C�HW�����'�AQgM"O�.�`N���(��\��D �+]~.�~w�_0ѯ|��d�`{��X
����aT�����Ɯ��
f��zG.�)5�oZgzW�3R�Yv����4-�#m����b@��\Ǖ|F�x
���v�=�l�?�H�NÈ>s;):$S��e�D��j�fO��\�D���@m��Y\GG�j6��JBL'AgMەW��emT��*�����t0 �i�����Ge�y/`֍�m��Pe+'�^Ǫa�{h�G��	!`[_6���%Z��@��N/�������-��kpGR��lU��`�n�lx�Z���/��W��*԰d;�μ��3(E"f�a������"Ff,>�E�a�o[�QصZ�.`���gF�	���qz����S��D>�#Яt�ݯ0=���U���j��o�M4Lg��@��☌�շ{5�=+*;�P�����9��o��K@i�Dl�rxNl����~uq~`��ZRM>Zc�L��9�ꅮ�0_�+��ܬ^�N������"��^C+��"��BEn�% �`�n���4X���YM\-!9]T�KF��?Q�D�j�.~#u��A# 䁴�\TrP�����RI�����`��2A.Dd�ΘCyN!*#,,�KKT6�3�w\���]�- gi��5"ՐW�Rk��o%j^!��6���������m�6�>�b�+���3Wj�l�@�۱�뭵?��^?� ,B��h���Q��tb~q3*��ٲ�
\�4&{��h���X)�H�t�JT�-u�h�$�����vt|~���ݹ�AWH91a�>n$��~�@\�����o��X�m"
��DſI+��}��;�aO��^x�`��U@?�I��ۧԚl��W���/7&h�Q��Lvzq�S�{�pZ�l�j9�]�)��zdSwQ��B(�	7R����":����W�*�	/��
��APS=�`)�P�Yl4]�cA�%�T��"���yZ���f���l�\j7�V��'�l��A���>���BZZ�A�0��K��w0SwC*P;��Lf;8��dMO�5DuzJXWx��~2��%1l ��~���=�b�(b��E�N���^�������PӏN�P�]�Θ]&�������#�k׮�r⮓π��c�$.~1���K�.�w�4p�#��O�f�l�Y��$�Q,��ɨ3�f��$�J?	��Ѩed��c8�]�k{{{���v=&�k�Ζ��?����>�p�T��J�/���;׃J��o{��� �Bd��լ�q�v1�Cd���Iim�J�6[�eY�<�Q<��-�b�N�}��s���аi����*&ƧP}����B2L�CI���ݺ�{��D�9! ��τD�����3E��	��fT�k�u����}WX���3RX6�'�H�~2�#������s�:���  KK����]��$.B�&�t`	��?l�8*PP�!D	=C1�S��t��D7���Vn�;)׽��"ĽeZ�<����>�����顐��^>��}��t�&� .mx���p���a�Lm�,iG6�F6j����;*����SJ�����' ���	��tU��o�b��˨'�/�m���k�>z���ն�U�]��Q���+!��f�C,ot<��{螘�G� ^� R;��@�n�yq
�
O�{�8}-��!����1C������fj��U�Ċ+q��-�����C�V�$`|�THxV���G_��h����V:�N)�ݲ��|��x>`�%��љ^�L�ӝ@/�<$ȍ5�҃`� QvȬ���5p�����y �9�VW�K\g��u��8]Xe��j^�o��S��@ǆ͟w�&�ο{����gZ�V34��Ds�6� z�;wrK����P_-��Rq>���p�b�२���R:��XQ�J���m�RQ������F����`Gb]B�����T>S{�Q��h��ÏpZ\0����R����L��O7��x��?}8�#�8�b�����N���C8�����D���c
��j܁���?u"���kѥ��.%<U:�/m$��y������o��?�M��<�ǠP���B��Tx2��蚘#���_d�RY�A=�� ��L���g�3L���}���T(_�t����~�5�����܈UJȈ�N��㶼rt���pSfXt�c��r5F�s��7~��~ ���j�4��Lf?V�##2���E���P�Ox渲ܴ��p��[���Rr?O�E@��S��Vߐ�sC[?BE|f��͖�a�^���_eA��Q��O5�o-]�z@�+IaB�X���.��n��Lo������(E��8��(ۍ��h�'��t�^LQ�e��'N��)q2b��C�ܟ�K���X�;+��디��M���>(�4�+��j�UtDP��6v$Q�l^���b�s�zo`���u��n�tJT�e �p����c��� �Fg���͍X@[�Ȇx�=<�y�l�3��.�^�b�9u2��K3���%��,���yc���ym�%NH|�(�+�ؙOB�,���x��:V6w��:��dc�LW��Hd�c���
Ԕ)�ho�G�IЭ���1�U��##�e�8�|������2lQ籨*�jX�ܦ�X�M��B�� <����{�N�9�Wو!�c�o����AF$�!~9��1�1!���vz3.e�4o���N�6���EPU�3x#�#�����cJ�	�rD�����S��E�$_���d�>���߉�3��k7�(��uэ��D��b�9�4?�*�:���d���! U���'��b̏����`���
�%d,--O�I9�5^�F���v�ޓH( ���o�>T�n�����TYZ����h;�32o�����aM�j���{�S���,�&��3{�p�%��� �l�����O͙�m�j���=�c�t����5�a=�,�Ļ27s$)@߉(����E��ag0.�@�������بc糬;ZX���mo�W%li�D.��s��[�C�Cݱ/�$�;ܳm�l�U����q`J����W��������UR�HC�Q����/�e+�}q<� �W��m�Q~N�U��X����P�9"*;^�Z�c���#��OU��6�ӨC*ܶ�N���¼l�f�2����6�; P��A�PC��`77�����%�@�L�IÖ��@ �z�ԡ�.�xk�M�c�Jm�K}X����CҀ�a�>���7~	��b%�q[��&�m����bv�F��;��vgq�&u�<��+�0�L�J� 9��e��i��o�C䨙�an�I��ڹX�.��:���E��N��,��6:A��'�k	96�9b�:>�ժ��g�8M;wX]B݄8����*gM����3��t|8_axLuR1��JbC~H<�Î[��S�&�=������7�I.��~E�M�O�Kҩ��qQ��C�m�Qi��_���]ѡ�i���#�`l���|�.����V�P"�3�̛�z��^7d� ���$ v�f�m�~�\W�~�e�3��]!�հ�]K#@U�U�>g��N͏�� �o��v�p$"m .��q#�76G���A�g6(_�l_�4�.X�֕��Nv]�JBuC���?�N0�^}+���V��9�ٗ��g�u1��oXO0A��W�s�?U0���(B�u(*%5U���&ԡOܢ����f���:�Z�A��u�C�(2��K��x+,�5�&�>�Z;�|L�X?0��_���U�v!F�X�\H���8.�qj��-�B�B9.�HZ��.tq��S�ڂv�k_���'�?;G[vĬ8d=��ܹ
c ���$w/��O�zN�>�l���y�LP��+BJV��ٶ���Hݎ���d洚��#��6�x��6�m���^����3��!v2��P��EW;�D侳�x[�x���9��)�j/=��h����'4�a4qy�-|��nk��ßSCO�3��1�8#q(Q���{��0�`��D�B�Q�^R�b'u�|md"�*�n��6���A1M@�O |�#AC�Ųݞ䫇�4U��{�_�ӧO��Z4h�Ȩ�ԉ���џ�I�t�ۇ'Z�uʉԞ!�b@���Η�������h$���O+%F�j��M��F�'q�D�F��򀗄��;Z��~���ܬ�: h��w��Ϳ#i:��F��5�F�+�u�j�,��ǌ�q�^<��	Gp��b����:Z�>j��C�S$#���q��>~�Y{���~����-�=��;w`y7څdo^{u����`fF�o��tbJ�Ψs�V?��R��R�Fi����yԞ�A!�)��%���E෡��"k����iw $���
�pd ����w{*	��+�<<w��^Β�Ld2�_�L��e���y�L�v�/�Y]��	˖�R ���hy+�m�J*�3ˎ�N��o��5콳�E��m\��:����K�7
�>V�6("�d� �J_�U)o^�f}��ia�.'�~��(�;w��91Y��ڧ팑c��6��T�-,���~ZV�|�h�9�F��S���D��*u7L�~���o�NI-�iP~I��B���G`�Xs�2���_w�x[CK���X*
?"A�#L��r��%S+�.@���@����+��M�<@aޠ���"�w�(v3�Өٙ�)��}�[.��$޳�3�
�tՀ��s%҉\�QK��T�4���U��d��TJE������X����Xq���:OA�q�A>#��a}'�����n�rN돎�5�7�S�t��K�`�����9yO�ׄsވ�`�)ٴt�q�lQ׮:��b��O4�m
9�������l�U�Aw�р*��t �����N���7`�Z����,�
NyO��u<���`f�۵��~��'d#�ws�w;<'�P�
��8�o����-�d�8��K������޽��������� .�/�ϘtTΆ1�Z���5Ң�,e����젎h ��>������(�p����F���zh��~t�i �"����������p�xU�����ml>DA`2�D0A��C��m�;���0ӯ��^كZ��W%��R����Z��OqOzZ�׿V�|�J\���Z���<�m�#�vK�?�N:8揎0kD�^�A*��!�%Q�?LN���{�1pN��.&� ��Y��j��,[L���B|��+S��Αu�d~y��1r,���z -	xdc��4L���H8�]�Ī(�&���k�m&�E�!K1���ذv�O���|?R�a\�x�l}jξ�;K�Xw�[�{�3툧�D�.?L5���������}���"����c*~j��r|C��E)9v����M�
����q��MmQ���[����!����ne-�������-��SAqea��站��<��ۙы�����P���4d\���_�ol<�y1Z�������b"�%]=�
وnƿ�K����x�Nf�u�~$�,3:���e�9�X:҄�{�J)��yC�z8�ͺ�K�XO�[=�^�������/2�;�:�D�1g��!Y��a�8<�j˿ՔM��Kxy��1m֋Ԋ����-���N%�'��S/�)������@�w�nǹA����sU��6L��6��~ԃ��m�/x��ۣ���@m�N��S���/U�����la,�'F1~5���nA�X����.Q�������{� �KA�U�sd��;�܅��@���xDM�q$�7o�*1��yᾛ�O��`bo��d�`s�I�ܥi�o���[��k{��]F7��,�g+&��?R�+���� ������� �A�X�a�7)&Ǯ,N���a5k�$<�6wu�q�3�3�����Vvz-�z��;�t�>���n�c�0ٴ��c'ԛ?�a�,��(�����G�tT�z�AB�ɸ���%L�'��R���%S���C�%�ǜ1�i�(���������6�����c��p����]@=>�Ÿ冲cE�T�Ie�7t�?(��0LEy���[#j��zN+k�K���[q'�MC(����?��������]�Y��Qx���S�j����<��p�梕9�f�� B� ���K���4.C� ؾ�	�2��{c&T^�{�kyaR(��'$]GW�)�)%Ȋ�C�d�`bY���c�$��}`�R,-��������Zv!?��^D/� ��-�r�ڣ���-��"���q���X|%j�.!H͂lzt��/je�o��400�����:$'GdU]ǯ�B��XS�:Z������"t�h�=��aqv��2�*x���3�Ti%�[��]
�z��UWn^^mfS�-֧��G;,WTT4m��;���S��sP����}D���
|���K�{_�s����X����2m��D��5�]B�)IѦU+c���l�B�U���	-%�G{J��}_�uݟ���u�;��:���<��x>�z��u�o�(v;쫌NH�s����A%0�x���)����t>Rń%0�B����	��������o�uvLo�����v@�����!b�]-�,9�6;����`��d�Js�n��k�u5%�e�3}W=fg��Jص�w*u���N�9�9�軿�x�@��� �k�,絳i�%VV�Y���=Qe#��0ծ�X���J�^�BG�|��ϯ�0�(ɛ]��>=1f�/0�d�V�G�gǕ�N��6Ɓ<V�}���p�,^�f��YM���Xcw�ga�Ի�=::t1Ci�j�y�cRX>:5զ�G����<�Hu���T	'D��8W�|sr$�Ư��bS$y"�P2���V,����f4<fG=�H
��-��m���T(ۄ݂#�����
K:ĚG<=g�'�V��a�6���� �F�s_x�['�wI�}m�8?�2^�+>`
��]�5t0嚖��sp ��_����%�q���j��N}�]O����0@o�h*,�9m^+�aA^��Gs'�� o߀�c�ܛ/\?Fȇ��o>YvZH������?��D��Z�����+ ��ڴ��BERI4�xP�)+�tù�9/���U�K����&�6ݭ3��d`݀E-?�@H�k�"������ةkiF�b�+��"�Q'�랞�=����d�[�(�[��U\�kT�ho?�}��}6�x�Q���?L��@���%aͿIMj}���p�����43.L��C�����>�h�-���RL'�i�����T�MӼ{�z]³E��5�v��2*
��@�)@̒��[X���֏�'y�F8�T��<8��=�)����hp�I��7
��]{n7�N�2�䊠#�`�bՇ|�,�5�k��lf�\���9�ۖ�sc=?��$-e4�H��e{����e6_
vj).��Df;�r:66�fo�lo��QtwEo�>���Gp	ƚ�i<���	�nEc[� ��a���S����7ÒKTE��xv�eَ�Z��
-�w�y���(���Lo�PZ�5�`����ɒ��%�-�#������-���c����J�d�'G������T`T��>o�u��I�Y�/?)cb��B;�VN�n���^��%=.�=�TC�����u�Bc
�w�D�.�������t	*A��PR��(=�;;M3�M��
����iV<x�߻���Y���	+�{,��2�϶���;l��k�.T�*��C/�tf2����8��[��GY�X��<rN�[�V �t�6�d4$xs�.�ݱs�\�85��м��DlĜ-X��ku��Ңb,}р����+�1���/O�����X^�M˗��}������~%U"�����8��!����[b��b�7w�ĐP�h�ƸNw����,sk���ak��s�-w����du1hg	0�$��)&En��W���Y�����]K�VaP��2�YЋ#�UL��<��l�p�O1��[���^�?Tpa�iRqHE���4+{���߇�]ad��]��O�����(0Eg��� �ws��?��H6��Ec�K���J�����p��.����.]��bq��e���w��X���{��b�
��S@Z�.r�o�n��m 8y�/ɍ?C�/ ����l*Bh��u�5�Sv����?/:GE$a���� ���JhT#,��]IQ�;�G���������-'U�`���c��PCׅ���d�'��/AF�
Y�F��\�q�3��v^�ӏ (g�
����^�zjR|{�Ý;=E��:=-~=�6�[6r�X�
�aAᩞ�t�;`K �G��g��*
�������n���ŏ��3��!-H�y.ͭ�\[:&���1�6����w�ӹٜɞbF���[�E��|��>1��g��5�L��Z�0��Gj&�4�P�N@�_Ϳ��?�s	�5�!����|�Zʳ��	G���O��Fv  f���R�^JII�u�V|�,�>,��������ʭ�u�A��LW����A��h)���?�}���ݗ;�N�����"\EY�����2�O��4Â�jT��$̑%_H���Ę+FK�o,����wqq�h�.�5GU��~�|�m��S��/�w���n苙L��~�?�ﵢ_�cX����j�`�#�S!�yE�#��1�>Ăn�h��U�ww����u��π[�r*�"�շ�a�]&�"�����Y������e�������o�
 =����Xה5XR\�h/��
'���: �R~�q����A3�D�L=וX�T
���_u6�N/�r�zޗ�q`� �yay%��)4��yHfN��+��"��n�$�jTѥ��M���4d����D�����2����n�l�6�>]��s� %
W�)-��w&����;g��ՍE�a�H��BP_/_�� )k� �n����������/SB`|�ܩF�R�1bDy�ݿ�鮫�o@�>˴�J�HW7�t�R��g���)���pv���^&IQ�J����̛�0���++W�֞=���T��YEĨ�8�P��٬s&Y�x%;� <��/\�1fk2�h>�ȹ�;S��*�>�:��~n�~nD���c�����*b�5�U�V\G���b�j��|�y�`fn^����J�y��aO��]��D�'�ݦ���(u���)0�
�F{��bf���\���D����R���K [�b��K��h�#��k�5Co��s����������؂�v�-^9̉����	����8���d/&��i��D	��Zc�;:hTvq)�`B���ue�����65�N�-�j���OƉ5)]޻��?���ij�'X4��'��F��a�����;C��w/�Rb���/G���>�ҳ����_1s^y=��9�ȁ�+��d�C8���qFs���h%����_Q����������4�6�<� E�@��K�ZOVc�̏R1����NRY�b^l8�H2f�Q� �fB�v�E0�]����F���G�	41Μ�*��~ z���{$i�y��Ɲ1E0�g�D�x�u
.+�IY@�rd��ځ�����gX��"��%+�Н9�ҍ��rr\i����(��kZ���p2z{��h�=X�$ɀ��[\��D�B�<<F4Y�b��r�P	��1v�6v�kLJ
����_䤝�M%�=P���cYN6��[3맅 SoB�-��8$d��6�����UQ�o��+i�GH�2 
���%2��e5i6�S�����[O�z�IQ��-��������F������Æ���y>$�Yc=��c�;��;d�tH��C��],OvI���~+�.o�`h
uE���4�'á,4���X����S�爋�ѷ�� /�F 0G���3�u��^|y㏠V�Y�Oi��4c�H)k�9^�;��|�͊�`f�- H6�RH��W� ��E�\��M��`|n��K��ɺ�?�I�5��O;�Dq�g��_[+{�P�54�l�}��ŵ5����mѶ�q		~$�*@�wV�!��j�!+�~��Ѱ�|v�6C'܆�����p�2CG��J�4Ao�ƽ-&�kƸ���u�?�)��w� �V�8�;s�n�#����@��M���ٕ�u@����#��i;w�,�&�ob�f�����$!��M�(V���֨)�j�ȥ{r��b�b�vh����ѫ��v�5�*��c�c  TA��L��Uű����"gZ��1^�/����ƣI���%C��<ͮ�ʏ����E���S5����B򅞙z��͇_�!w`��b�#�4y����B��AAAԨ'����9�f^:��@���h���_qS�Z�[�1N�1�AB�Qh���)=��
��W�}�Ġ������F������2胎ֻX!j 	�>�D��ִvW�e;���s�Fr���#p=Iʹ��X���߹w�0��ޗǩ���w���t����L͑UG\̦�����Ȫu�#@ʘ���`�:�
/�jnf&R�����ո�{����v�f9IP�Bө:�4s��]��z8��
,WA �[.|����diV���"�xkt�s�u� ���i�k8���ze�:	]/�(�K]Ĺ!��p�zna�Y<�ӌ�1A ��B���/�o311ѕ��
��ɿ�]8=� �w��c2HH�4�� ��}�A��Z�%,���:s�(�Ȋǭ����f��	�ˬ�]6x�h�����P@�J�h�g�1 �����.��$�HU���߯�����,8�����\V;9�͇�j@Q�0���BT��w���D�.Rq�lj(R��4��������p��{ ����k�����D�
:�96����#���&J2�4ﶶ��7*`��i>9�(�s�)`�&q&�r��+z5n�Z�n���o.�������=�kb��ps�&q8�W�8�����x�(�Bȭ��]�����U"R���;@�|G�ʇm���T���Xh8����U�!�X"�a�'%q�7��G�{�������s3-�C�Nz�����VJ'�����~�,emG���@*!A�ZE۬=F�LXqN:�Y��c!2HOD��c�&k��	������*��e����.>���	M,�G���+�fU��C��M]�j�N�>e��_�͉��0o��n�0ֈ2�ѥ��v�D�w^��؁�`��ڴl��z�SÔ1��.�4SS���ڬ��>�X�GK��@�ڵ��#>2����@�t�X��) > �m^]�����$�L�q� ;^?Sϸ��&�hk��bx���8�v�\�����	=��$ʋ�>�d8����$�R�FRJ.	|�a�:�ũ��:ߓb5��<�o�ϐ��@9���@�T�C�)��v�I�?r��7�9�{�m�sㅅ$��{��z�"�&Y�\E����_����G�N��Z��L�߹�tUq�#Mjj^�2�C�Ejr؜��.��zk��:�eO�MC4(���͟i
@̄bRq�&�.���&X�F���ن�q�xX4��g�#��bf�t���.֑7Z�)�쓔iɃ��Q%���saL� )b�^SPdl��4��U���
Lҏ��;�gW���W;k��]��C��f-5�R�Mox�ڪ*^�lsް��";b���ܢ�B�n�������*^�o@p����k�LP��^%%%R��>j�v`��&hR�CM�qE˹pP��4����2�ۚdj��E~*EjZ&14��Yg3������%oT�kIi-[�y��
�|������ϋ(���))$��E�ԧ��c_t	C?f��9���$Ji�&E/)Q
㻓�O���Xl�{a�ʹ +"I?V@������&�N4�|�O�.�A��@ ���IrR����D�^꤂A*� ���(^��T~X�|#D��:��L��rD�U%�`[)�$�0g�諽<R�a��`��M�������mF=���r;Ek*;�:ͦ9IBԀ$2=$���Ø��ν'�P�X�<}�zIp	��$��0��S7qyψ
�~�
��D� ���}XՈ�G���Z��{a�'��fVV~��НY�����(��e|M�nx�.t;��)X���@6�v���9K�Hp�J�{����J�U�:Ds���(/��̣�	w�o�־3�QThYm����GMR��#���Qdm��;	$�s���_(X�z�X3��dz[0B��Dm7���Q��H��}^��,P��od��"F�{�5C��@$C�(ap�}I� W�vJ�U��&�} �ۜe+c�7��P �H���Z��h\�1s�N��5�f����朱&r��/��*��Q]��JL��/~�>A��̇1 ����@w=;���$����a��:H�gz�P��߇Z���,�*�$+�ڈմ���)6,������D��O��'*v���A��N0�w��׺_� �K�`5�*-ޯ��o��l$כ�.���=��
U".}���}ٲeT�a8TUM}e����̮$�h�`D������;�UЉ��Ō>eZF-tl��G��OG5ͽ����.0>�z�J�#4��T��������1.6�K�Q'���a#O��ы�����tĳJLL����ğ/�K�sz� � ��}��M�v�����vf]��*yg�����1}�t��Km�<�(��A\��F��,-�H2���>}:�]�"���L{�ɾ�?���忘Qn�Ҹ��NH�Y���,�U��t�-����*5�E8��vw�:�?$�`�-+�DQ�B�⊁�!I�\��$�>�n�tޢīV�AT.$}�����??�|y}�`Ѩ NC���)�I%{��m�	�U{{8l K���o� .���b�G|�/vZPU�+&}�		��?��m%]K�9L�~R�b��� ���R�X�O����dT'�}��bi�+7������$��X�^H�Xk�,��H��R�V���M����������L�ъ�0,���^��U`J5����FL��R��Q�a=��N?���N�oO!0��� ����-@pr&}6Q�#vӣ�x`$uv�)k0���� Zؖd��d�H�<���ݔ@��Lğp-J/��B~;aR�q����+���I�oٜl��g�ja����ߔ���Gн�>qi�M}6$�?�;�Zj��1��\Q��k�9 �/I9s��&U�+�coM�fh��^d��Dl�����f��ڍi�g�4�E�4w��F0�����Ԍ_��T���L��8C�M2.˃FB�}�}����gb�ňTa1x����������5w�EH��R����\⴩��~'�Ay��Wz�&�d?Au�����ƴ�xP�x��:��iJ���������X��JJT6�F�fn%��/���؈�t�4�~|,\����ǊL���Γ�P��?��c�Y��5���;bb��s/����?]x9��_�:ijw�X�_�5_�d���>w+x��Hf�5B.!@�ҿ0[�d�
�ӓW�,�+�<�]�p�%(��;�f=)��~ɫ��`��/�Sy�ޯ �aA8�7IM�n	a��0�k�^]a�T�J��#��D@�	n�ձ8�G늆��NR�.#���,q�r\ϭ�s�";O���� ��k&��N�����a�+��,�d��e�Iu�qS�?���ڀ��Ɇ���g���%� �T�`�!�T.�:�n� l�4�-��е�
��OO�t�)�<��ĊV�Bq���F��f݉YDL��痗0s�ki�Ϡ��y9�8�`�6��no��|r����c'ô�n��u�q��2�eZ�H]��k���N���8��Zj�H��Aatd�*��;@���5�V����I^^+���R�{�	�Q�bt���Q	�V��� V����V������ټ������k+���������b�6������a���AT��LUTBBB�c�pq�4���%�J�T?<ʸ�B�+
A���k����$ \��o���:���0Y�?�1[Lv]��cݭ �q���A� �aʝ��0�@RaR��1IA�"��NX߇�0X3;��I׿�0f�5	�ϓ��%�	~���c��T�NY�c/�C���W��N�Ǯ@SW�����)O�h��hc�j)�=��Eʽ����z���6�Kk�T�|||�x�-K��+1</@.!�h:	�JCJU�"��E�f�� �8��m���40Q��7!���1��S�ͯo�cҔ<y���]M��U��Yk[*O.�~����m�M�Ci�&9��$b��xGK�2�B$%%�B�� �r:�(�� �3z_�eJ��yI�|�M�C���������m��L�Qe�6�Y%�i�&p�@�N�LP��V��)�)g��"J(��666�p����^	��YY�nkJ���
}x��%�n��C_�[3�jk�a������134}�?w�	ӝ�Į�n`����`�ПEC�<��gB������x:I�F�)%��Y8_Q�@:i�tŰ�����|.3��9�8��̙��A��NI���C�-�gε����4��r>��y������l,��w41}�7X�4�܄Gp�k����]�[�"�W`tj���!([A�
�(�������!DXwjCp��J;bF
�`�l��8�9����%��XW���^@���\0�!��߮�o�œZ��:����с�o�oT�w���a�A��ra��𾎩ƑA�
�D���9��3mjS�=��ȿ��%�⽚>>~?KP��31�mn�����Q N���4����t�Lue�﫱	92��*1c��/�k-'�}~��_1ƴt��-x���ԛO�?D��&8�O���}�<���wfH]�6x6�I���Ys�y���?�9�e�w��9�Al��
�~�2}ss=}'�%�U8?7{)�A��)�PM�I�,3|e{^�R��*�=�!�vG� d`��^�cv�J��G��5@������88��rAGڗck�z��;%77�ٲV�,^�`t�gA[��;�Fp�`�A7b����&�;U�8��Q%��+�y^"�T|�@ Չ��7/�Boo�I|��G|f�F�i)/>�Z/��FyѢ//�V�Jje��'����\����s�7��n�1�4�h�x�}xo�m�GS��N5���s�(�߼?kWj���_Υ��K��V���������{0;tމ-d�VMM�D����2a_o֦FDl��VR~��a�
��'JH���	_p�����X>�TZ s�.��j�����/@���.~��̋�7(ʌ!�0;�]0��Q�J%�F-�	l�r��O'��GGDDD�����׬�i^F��Y��kD�6���c�J��M�U����-�� �[-�l���~�%�s�a�wL^�C_�u�l=�R�ǡ'U�L��\-%%�uS��]^���گDj��o��/���vy��x�̦����ێ 򳅮�d�LO���?����?�f�Ut����"`A7�ď&��	P�FW�U�PA��FԦDGG_ś@D4���&8-��"3/������Ǥ�~C������VWWk28�w�Ύ�)N�!l���]
!~ڱ��aW��F��	�ˀ�&c4;D�D���r���: ���%�����fj���W=�]�f>���NJ&D�AQ����R��F	��nJ|�:wơ����������1Sz�\|i����Ҥ���ZX��ط������kl���7�䝊4�f��x���m�Dh���t��p4>��tl`һ�­�`���*��g��	����oa[�;b
Fi���;�؁�����}7H�f���=747�9�0ݮ/�x6ô����1�Th��76�X�8�Gs��W�7�F�Op�wE|�o�x'SL�
�Q�Gk����S͂�%l����L׏�H���+;L�XfƝ�����v��3�}��捕?b����w�����=uJ�~A��@���_9H��&��J<A�27�J~���ÞaA����`~�4y�3/`N�`��X5��s�wK�hs�H'���{�K��-[���Q��x��R;t�X95��;
�U2>�֌�H�
#�ќ�1��������ӛO:�wjm<�W�/}���}�zL�jE���@���mX�/õ�]� ��k0����O�'���~�8�!�_s�Q���,��<¢��A7��Iw�����Ԫ[r'�-�ކ(���*��}�� ���Z�:A���+�u��d��J$ɽ
!j�C��f�j���� 4��E�{��{���-�L�I/��DV�)ǒ�YS��z]��̭�����ӯ���ZB_"#�n�AaV�>�}H;��ЧJT�����1�a{>���������7���|Wt;�%�7���2���&ø��%f���Xd��7�`nU�3/�m��`Gg>=��Z8G~{�����8��5&�FQ+!��;�ϙ"��� ���#�bW���r2��Z��}Eh]��paz�#e�7"D�2�/HaR�C��D����xx<i��iџ�B~�HK?2o���/鉝Ɨ\���L�An<A10��0;^�*�DM�����c��z��_�zj���??a��X�j�偣>h&�f��t(����;�
��������c��=���K���?�`Dn���J�z3oTY�sM�qU��7c�����#���x�{<��������~/E��<�y�a��2�ߌ!���덄�ob�>�<��Q�^��<C2��Uy�&'Km6Ⱥ+�{���0������L���;�v=��<�g��������X��i�) ����,�ۆ�}���Bǰ�w=�Q�֫��L�?�1���$#}�\l�����������%�F���-Rъ�JFK�_[�hjy�nJ?mFY�|i^��g��1y+�m>Ǝoզ��LbQ'tT���9�p�|�ҥ�U�zv(HW�L��ȧjA2R'K������C�ŗ���=E�s?�!�L��ʑ,�ڳ:$a� zh2�/��̴����񫊊Jo�=p>�=���Te��s�pz�un=�~<P���&f ���>VF!$�0��Rt=۪|d��Y�vu��N|^����!�d�ôq��K�k������0r�r�U�����ʹ(z(��+����cl�lB��=�C�VHS��l\��n�Up
N�+�
;�V�L���o�	5����"�p��X�4���$�	�tU������8�7��/�����t^�G$����~9�N�'e��o��-5��WTTDm��p��"K"���+�m�8�8.�7�\�U�*B�41a�`�?��1o�<|�Bd���O��U�8l���
a���TЭ�yn���+���g��k_�R���*
���[w��zKuM%��w�pRY��p����ş���3{��b���Q�ZB��X�w�]�g���p.����
ȫ�OS��k)u�o���cN�ܒ������������W"`���= 2$EhBj��~�} �����CRR�H�
��Yqm��`~Z�W�Wo��	C���w_�	�LLZ���`���1����mƃ���'i���Z^�k^b�ׯ��6���OL��?2yȄD��KKz�LA�
�P�7<<m+z~�/cw���p�^|iJ{0n53zeS��UR$1[�7�Y�p�]=�cP�����h$)Ju�L�}�7����L�p�ߴ�=��V9��_۷��ֶ���&���NL���,!i���D��Lw6GG+�p�5H|�8���qG�6�rN��	jf��Joo0�O�>}�Qp ��ŇA�q�z�"P��a|�)�w�������z�H�0�b �7-gWH[� I���]64̰��3��z,g������K!V?�� l|�~�ky��P���٨i�t=a�;�U+���o��n�pd~z�!ز�>|ϵ#����3��&�L���Ejd�zR��TYY��9©u�X�ZVV�`�n{o�ZP�8�鱎�j��*�OE� �l,��p'��D���5@�}��+f6kFrU�띊3͊�-� \�.N�[%����5S�%���QaM#5V~��H��!B)�8�&��C���=Ht~́�WQ�V�፫���mx%�/A/X�@3���^[�g3o����@��PaY�������in�I�	�
j�cυ1��E�]�a�6???I3�Y��'))��5Vo�k&��F?s���"��/?�j2�SWV^�)q��_A���LK}/_�l8nk��U/e�oƨ�.I�|��v
}����UO��=z3�-8 (//U��E�d]�o�m[h��ۺ�W����E�����1!��6�9���.��E*Ʉ���|�i��O���5fziֿ�+
�z�h�u'�>%"�� ��B`4��+�������7�B��#��>�ٷA��B��=~3�|�զ�m4_,!�&��t��Gz8f]�M��׊u�5q���I�?�G�~ML�/f�\�~aYe劺�:�6nw�:��Dp�W�N�(m�\�]�����ש�О�ύ(l�ٝ�ĕ����X��s#�FF"T(z�������U!�� V��oEEH~�R�k�W�Z����N�M�S��f0�l@�wv^���i���ъT՟}����'<�V��Y���a����A��qw�w��L���i�'�|i/����D��(ni���vM�q�`t��%a4T��-_���9�%�K@��V��ǿ�BJ� ��ޓ���z3��@��ں�>#u��{����#�˛]^�|{w��DȞ��}��$>�$��FS�_��*Jݪߕ;7.=��a�acQ�!��e��N��V��J�d���_����E�~{�P6�HĪ�
]�EL�����}�B��$aQ����d�����\�(��}��gO8�`�pҹJssw"�,S�TQ!�׳�s�A�"��>ԇ�ǎ[{���I�+��5�-�K�Q���`g�`ׁ7p*�d�*�sڂPD2�љ���"�3������[�� ����*���ӕe�?��bs�ͧ��6���7�h\�������=���_Ǚ
v��Y�eL0��zV
��鞘U-�ĩ���v ݧ-Ÿ���3�k�㏽9����jD��<���@c��{�_:��Gl䩛��Ӝ���$��0NN�+��!�B���eT�'臏�c_2�O�Q4����Rs�_a�c�E���l�O~,��Ϝ��w⌋�#5�����Ok֮�{'���f��짮U�ߴ���r��l8���Y_�|�,���i>uqA��#�,��X!�f�:J��WPQ@<g��ʨ��Y���~!�!L��ǀ�B[��P6x={���T�6����(;g��6�Ź	�ш)P�Pc��?D}��j	�%#0bg|�wͅ$#���p�(㙄����P�aأ;��,�|�'�<פ*�ƘP��؝��M�qףd@]�/��[��2?5������I	/�:���A"A�H ���`a~
�\���.F�L�<��ŅL���Z�փ$i�&cpmP�U�`ۋ����q{e�*p��6�������ͽ���}[�SӢf��Gd7��T�2"�s��bY��)�w*�������ǻw���qI"����^o�)FP�ŋN_#��V[�!do��$�.���Y�1\����I�����an�����Ltx�|���!߂9ɕ�X��Sya�B0-��`���=�����G�y��%�.&rc�� 5�����SV�"=ommeNK��@j�����h-���֟w!e��Z!�"V]�Bd�m�vV�wuyc>n��a�K~x�ٴ�`� ,��[Lv�D=^�wW'��Y��	�*�ӹA��i� �ga!ݰb�%t���iҴ���foX���>4�"K�_I����c����>��a�t�����hT	�>��_)*��o}}=���@j�-��A���
~�)�����r�T�,e��ѽ��E�'6�!�~o�k�yl�`łL,Ȳsp�(�!�����/������xˇO��#+�Y�h�b���`*z�u����$2�ϔc@��0�˰Ot�Ǐ⨣D�{��F����0�@%uw�~���EI��h������u��={��̿'a:'H�Ѽ0̋[� M ��T94_�8�X?u���pU���o$:���3�X��������ZB?��,�?^�!��U�W{�#�<E)�һ6��AR��������b�4C���z�j�����}q8��`���à4�0��9-�ĵ��x,��H
�nC7�%��Z�<���L�ʆ�.ED��	�Z�ti޳R��LUgN�Ɲ�;���D�:uꯠ]Y#է1��.��1H%?6.������_-�����F�+��ԘFVYE���J٧O���rPA�-���x(0�P`����1��ѱ�P<SL�����
ڶ�� 
����`����Qc�8&������B�ۀ6	j�H���Y�;L�`6�2�;�G�ӱl��L�cӈO��g�����rr���@��J������ѩ�Q2ߛEm���)ժ!�5����@$w�L@\!�q�o����]��򮇿$�L�c-���0��;����wj���Ԭ�d����*!:������Bh�c�����R��̦;��o��ݰ���;���k���RS��?�*U��x�Ԃ��Ʈr
�)�,��1&�����28�ڷ��'�� ��7�R�0|�]�r�����&?�(�t�6{5>�f8:���^*���K[I�5 'O8�|��u�믉�%y���24]�<�(��3�u� ����� ���k1��ly*s�/���G꺈��q��s�����q֧�OY��>e}��������)vU'�_r�xt�u	����;˃�b�X�����mb��w���j�Z���j�Z���j�Z���j�Ok�}���q]5c%*9b�?߇�X-V��b�X-V��b�X-V��b�X-V��b����2�����o3/V��b�~�t؈���y��׺o�x��X-V��b�X-V��b�X-V��b�X-V��b�X-V�rk�C7yL��uڰ���5���8Y-V��b�X-V��b�X-V��
����w� �m��j�Z���j�Z����J<]HЉ/N�E&�m����+�;~�)��j�Z���j�Z���j�Z���j�Z���j��lї������~_½5��Ĺ�������c.Z��׿.����;��)jm������������������b��5�����>~��?|��Y�d��5 k@ր�Y�d��5����kzz���م��5��*�ږ�Kt|��k��<�f?��+ެ���!��.N��]k����94���[}�缸(�ߒ�����������Xqa卤���lO�iK�y�+)Ŕ�Y�+gP�}z���g�{���I:�mZ02�E����u�.��f%ۧ�E�GJ��&KO�5~�a��I����O��Jac�0�۞�O�^F򎰓Om�έ�GW��|v~.s��ۤ0���r��&!8��z��:���-EI����coO��9���c�.r�8E�����e�ů?Q-��x9�����E�F�=��>s��&^"�����cs�������:�\�����l��u���x�H[k��F�f�V/N؋VT�z����1��_���X�7��0/�͉3=חYԴ�2���D��X�����j�������lΪ<X��8r����6_��r戡ai��O��ZTӂ�lmm_�)��w��,�z��tS�y.����̝��q�ec�=OՌ�o��>?�����N|�t�����%��$�a:�t��ٸy��~����>7�_���HW7�k�� M�;ǂg;>�R�Т��7�ו��46����̭8y�^�/�%i�Iod�@~�-�W��E�5nc�M��$o�Rt+�u�l��i�A����jV��:g�K|9V$�m��� R?~l�L�.��/��;�� �o���F�;g6��-�ӧ�'>~�������
�m��)�[��L�2�~�&==]&\�A���'=!>�U���Gt���yڸ�٣�����׀p���Όq��J#:3�;���ڿ}!,�f�y�\'�VK?����t>�a��3�ڕ��W�mH�5��[J��Ţ���O~�ٕ�
[��G�pv
�	�͖z�t���$�ky������b��}ʀ�{��v�G:�6���_��^�{�d��B��7)�m^����f?E����k)�ms<�olf&R�(��I7۫�*��x]m|H����N�뺉6����]/^��Ñ��Φ���،tU�Kv������K�����2��.J�x������	�T�Ġf_�G�^�G�3�}ԙq�������\ⴹE��k��+3kA�]/�P�V��Z����@��>����^J�nW�|���xk�ۄ�YSa7�>}S+9+�E=7#�]��	U?�[��;�u�6��{�+2��c^����;�-řF��11��H��;��J��QHk^���3#ͩ�Hn�=̦�6���nq�|F��p
͵�6C_��9֥ɇW�t��ON���4�O�q��N����}��6����@S�j:v�����+��efw�E�B�#l-�Ͼt	F�i?M�����fI8�kz������4ڞ����NjKuixCo!t�����ʫ�Gw9$�e�?��Q���o�Ro�dKB&��o�O�N�iJ���q��)zy�O�>m�y��ѫ�=,��,}��k���V���A�Ӎ��w�5���� ���କ��=fݍ��sMlF|s�-1��T�6ǒ��.�9��!��_Djɒ%�[����t�4Z�^�8��у**ð��IfJ��;zG'���
>b�O�n}zbRүbbbt{��c�k��-GYK4,����N�h������`[�Ao�#a#777zNK�e�ԇ�6_?��;'Z5�|J�2�1�jp�2F8���Mv8�^ͻZ�k/Gyy���	w���������Gdm,��T|#1���mw��}��;&��{�;̓��T@֯2�%''��p�wg_,
1��IIK{�x#�������Z%SSS��Zm�jj�������V���ݹȴZZZ0�����t̳_$��d��d�}a���Z���=���L+�k��G���?�`r4G�� ��ɑ�k��çj�)���4!�6g����F��2������8{5�󄄄��`���c���읾5�ւ/\�~hܓ����C��D|S���O��*�}��mm>4�T�L�>yy~��V�ϴ���oLA}KS��IB��o��j��WY�h��t��u@'��`�l�!ضQAQqv,ѸP���pL,M4&ԧ_����w�;�LL�>|xmӁ���4��/���6iUf�ո/ق/�L�U��_�:�[Z�,��u��o٧j����S
���1j�qۺ��Y�&��e�5�i� �<i�q���w��i�O��b��;�C�u��I��*�>*y>]k2�u�BBf��_}nx�lYm[[��sק�%��n��O���+�׺�u�#�`�wZ��y$����kv�f��#_36wd���I�ګOO�A��m�l���	ǵ/5��'w�^ �P�J_ۤO���)����͈�^AW�K�b&G?.&�g����C��S���x�Og��K��<���C�}��˫���W�g�ߢ��i��>�笞>}6I�k��t���>�L�������'���t�G�11��\h5>Y���m:��^%�c�jI{��:�[%&�2���c��;�7P�w���i�3�:~��#bbr���{
bm'�sN��q�
l-��ˑ8�86�Sth	�s]�p.�������e��b^F��}�˛��5�<	��Z%[�P�����G�6��}���c��=��r�Z�M�Kݥ@Z����-��
F<I�*�5�'�j���0[	�I��I��0���t+L��=��w���q{�/<�Y�jn��I������P�\��g��ٔ�ՠ�穕kV��r�2{����I�^�,�֞n��F�[��3�E�t5�Z�ͼ���N��/>�{t
�J�)����Ŷ��������I��2��O�4����Z�Lw�I_�*��76f�;�:�a��(�zy[��#T�g��~�v���h,��S�V��{ԇ�N>�7Շf���wG�Z�r��_cl��,CD�#��	�F���5���(\|v0o$�#aw�bq �.��!ɛ���tw�O���m0���E���������ޙ�gާtG���+V��EŖ�rӲ
��ތ����:��=5���d�nS��&]5�V���j�=�9p�[�-�� ��vg�x�4���ڷ�@iK	}�߱x��d/�#�3��ʄ�l���"�C��Go��JKJJ6����4�s�5������XT�����bZ,RŜ��=u���+��G>�~ASfC� Z��ԔU���8�9�~�T`+�Z�B��L����RP�ڕ�J{��N3�e<0bG�ӧ}��̒փ�'���"�B1k��Տ���#����&�<5�q~}z�e�0s^w��������&ؖs)g�;*��3�g��3��M�}];�ӳ)h�䞨N���>ڻ�%,bn�pB�"�Bސ͈�ğ����tv�ff%�)*�g%[�m_�#D�M���i�Spnɽ0/zc1�j8y�XV	O�X|�<RͰ��v0�(s�+��C���5�n������ӛb���%�ҵGN����s��@`��-�0l���ƭ�%R*����g�t�C��D&����m�>�e��צ�2�&6u��W��O��.�4|���qd���>�6�~7��\�S�3����Z�"�����|���ۧJ��hv穔<�1�?o��$�:�ڹ����4
�x���7G��i&��g��ݛtɮϖ=��=E�;���05��@6�K�E���RD�q6۲c� ��Y:���R�w�?���t����8k׭=y���᣷#�������G�f�R�j~���H���HM�R{�ܾ�,}�cǜ��c��}-�iv�q����ܻD���u��n=��uqo�^���)~vN(�b.-w��rI+��Wzߑ���3�x���k
��͢u.��!��^v�ҥK��@����ގ����T��}=�I�#�;'F}j~����?��y7(�m�ל��_k71���/l!���wH�]��լ�<=���	�GT���~���#G�d	)e�nDRb�z��j�H�w?�.�l�I���l?��m�[���I�=Rк�"�F&3�u\Nh ���'`�U�/0ia�����h�mi�#�z=�K7�6h�r�$ׇy��uh {�}�gdZ��^fg|f������L��������Sͭ�v�I���p�Z{����vC@�O�vdXrqH �ؒN
`:���5�96ԉ����2�ҮN��]688(Dּ�{<W~mSW�3׶ Ǐ`�߷MeΦk�EM|��l�ӧ�rH���A�lܴi��yĊT8>3���m-j*�N�4�yl#_Tn0�_KQѺ1����X�#a�h��5)j+��{�Њ����8��B�����QP��{��ro�����0���x�&�N%���,�	mN�8�m77�Y.�a����/7�>���Y�V��^�#�[,�}PpT��6��;�?�U��6��bY3{?b��o�Y�(�����Wi @�q�Y�,��m83p�þ\���^z�;D.e��*��rX{��ޞ�qg�����}��:�~\ץ�w�����-�)�-|uv�[@��\z\��=L&��N�Љ��p�`L�m�1���g�,��mrt��og�8�,G�v�C��ԏ����P�:�d�J���ه��0m+�z}�]E&��@8��-a�������W�tF�k�񖜣�v����g�� * Cq��h�#Ge�^��-��Ϯ!+=��P�U`P�<� P��y��-���v��(V-H&9��xl�Uԉ]]ghf����.h�;w<�`oГ-&��q���I���n�n����壷�{����	.y:M�}�����mHWϞ=7�i���P�Fi%7w�2��7&/î8�h�<�S~9�)���q׮]�N~��=����WWz����b:�~�:~�*t���ם&���2X0M1|��X�x����L�r]�&�Ӣf���˗V-��o�s~���Gh|�nP[���S�� #�U�uNՂ��ګ*F��N�w�0O����s39��,ԙ����\���^�=o��YM�`��d��:��w���#��i ��Ig%�=�+�	L�՘:�@ϔwd�ݧ�����:��E��&}D��':����6�17�-U��)�5ܰ�w��=�Ik��:�+��}����������4��֮mAR�^Г����:+��ڈsv�7�lG5���s8��ҲG�G x������CJ�1�I{�-�;2#^4V�j���B��%�nKV+������~P���W�ק[-�T�Y���wc�}̫+�L�Xԏޞ�����N�r=��{�����{�b��6�Ӌ�a��:0��G���.�B���엫�B�Adk4yӬ�/.d_>1=� ��Zq��/s���O��TVL��	!�pPf�h���]����v��7r���P�tn�ZH8�k����w[�;+�u��-�6+@�uD@!�G�*��[�K�>���T<�#D�q���'�g�߾{��,�\K��ಮ�.��x5�u���ޚS�cgA� 3ܴ�|E���8rğ����>7�����0'���m}zĴY�RG��=!�i2��Q��I��;.��M���z���ɲ.{kRN[Ը?�wf�]$t��:�� �����vefL̄)��~�4�Kwdl;Ƣ����(�s�:��
�6L8��?��q�Omm��sC��,��w�c{�/$ކ_5��ޖ�)5pq(��rF[�b�<�!D�!*��fE��A0+�E�����ή��0+��5���ka~h��bX�������e�`��l��+?do�9(QQ��n�����q�Ӟ��ys�9�6|2!�k[����)s�ɷ��S�n��W���]��OI�yl���M��ʙ����e�v�M����v�����y"�o�)о�J`z�~�+��E�ne�k�Lм�)�v�����b��3?��3��"ϝ�3n޼iL�^/ϦF�[�j��"sh�>���.����wM�\z?:2�����~k��&Єג;�������	���8P�������i�b�6O�^{{�� ��S.����ۧ���N,�?��i��D��4���v��?ƺ�٥sz?0j�-���r�~�����]�~wO��~k��|u�y*���>m�zfkZU_9m}_�z�ӟ\S#���}�L�uS`��C��K����t
�O���+'>8�[}��B����}4�F���^�c09�EN�ܪ|ߖ�{䕹��.u�G���I���{��3�%6�w�Kk9�T���^_���������{:��������^<=|�4]���ze��iͥŮ�5�K��ܖ+����~��݋�A��N�;'��ʾ�ǖoy�k��)qB���S�
~\�H#�_�n���}3�No�������}U�+-qu᪟u���]�����c��9���e��ү���z]I?W^���d�9`�;�H��v��f`�ڟ���J���?�_�SjYn)�(OW?�uN	M PK   �zxXp+��  y4  /   images/f9f29454-e4d8-4baa-8657-cb66eaf7dadc.png�{TSW��7�R+-G^��Xk3H5 Btԡ�mu�!b��	�5$�ڑ��UV!�NeZ�GyJ�C 
H|	p �B�ȃ���}����ܵ�.X����w��������܇;�^u} ����0`v�+s��ߧ����}�gP���~��޸c# �����9����?�`u�k�Χ{� ��u���'#T=V�w�CZb����W��T\*����z�	��V2�U���!�����/ٍ��������âd�C���z���?����C_��+2��sX<�:��3\�Y8p1z��X�%�ߖ�`��+b�j�p ni���͸��.mc=lX0c�1͘fL3�ӌi�4c����y#�����c�>)Hr�?��l������yXE��Ӛ Ir������0�����eX- �㪃��Gb'�YV�:���Q�4*�ˎ
��������ŴJ%K;�k�ʰ��"�����|�Z�=t����t��,/a�b�rD�U՚��D�D�xR�mwAg���NF̝���X���g�h1��A�H�������}�ߦ���R��|��?Ǌ��ʏ��V��]#4g��d ,@B�e�/F�'��)�\��=�F���3��������[e'}�5�#�Ũ1���DEa��@q#e�k�ĭM;�@�6<p^^�~Rb���9R�������,a;�����ȴ��B�������ܴ�}#ny���HIr�Tm�G[O_�
Q�n��U����|���T7Zک�IyՉ���%����`��dTz��Ȟ��e�[�̓4���}�MW �8#�CZ�yU��O��Z�7��B�Wa�#�ܹ���H�ߦM~��*�p����nO=�0�Y�*xz���M�b�ތƑbi9߬/�|�?6 �X:�-S���'�X����Wc\s-#�w��:�O�3�5�ٯJ�ӛe����ҫ�	H0�1g�''=h�&V�_�o�#"U��Pb�kt

�7|��I�x�)ω����4v�'j��h�xt�Y���~�D�tw��)�Ni����W�:P�mM2sQk��)�~�B`_wI��� ��44`K��|F�&�ƿ�PWcT:�?���Fī�������˫&�K����OlA�w�^m7�Ɂ�#��	%����6�8I�	�ރvYn��GZ}o�IT:;#���cZ]��7���:ݹd�ii[�h�婳�]k��Q;�X�o�y��U��^C-��u9�|�n��+���MRfǀaR���@��	١�(Z�'�h�[q��h���6�7j�p+�9=|��ugoo�mF�#j"�����Ջ
O6hj�|�vg����Ll(r߳�(��;�5���P�XS���9f���Ugm�&���F*��Mj[��`���?�"0J(i[���U�M��/<ޜS��o�rx�.�t1�x����X/����M�X�G@�����1�ɬF6�j 8r�S<p�?�d�~���'���%������QeV=��.���θ����иyj2Ј��h�]�G�mL��9����]ѽ���.��M�೨e���7w�΄�����6��Ȋg����CSϋ���=䍪�;%xH,߳��%&8��]Ζ�*m��l�N�i��>��kJ˾��sq-NQe��qX=r?��� x'2��!�T.~9��v�Ԩ����p���3�����}z��yz��� ���	�ޝ��2�9��o��~=���P*0��wY�{�ϴ��p��=X`��҂&�H�J_��PrYg3�8�������R9��B��*��[���Q^)!_/W���<�.MC"��d�p���Trg�Ҋ��G[���8`>�'�6� ���{'����q��6�P[#����j�
)�5b��cy�0����1`�_�d��^VN��?agM��ژn�C�T*�ҋ�d���v`�?����L����p��0O/
"��)����!RO������t�lz���[Le1>�������(	f��R��S�1+�����#Ѓ�c0u�:%�b����{�?\��h���Bs�;,�X�|a��lǽ��?Q�
:��a�l�����i��eD�8��r��7j�W�;��K���e�g��k��u��+���!�E�}}��S`�Ҧ0��r�a��|�������+b�"W��ܑZ�Y�=1yM׽
��5�;a�g��7R9	,?2�E+@~���h�EؕV�,�U,*W��<��W�5OU��7��D��!�V�G.�w�&�m�R��Ј5����A��m����A� �����@�������'��!�5[Wb&�$����O�
N�x𢝂��t1SCm)���R�0�/?R�@����A����v�ųNH��~�ƾ�p(PmR�g�q�v�*P˙2��r�� ��1��"+awY4<��Z�p��a�z��'eb莓in�j��W�Ķ7�y���ꗀ�[y-߶������wYK�z̹�0����*y��o"�XZ�]���v������|}�ȭ5�p_"#FdCs��t#�+G:�\F_p�R�a��9YL�Y�����zl�񁋲%w�"�=������'����j!�A�d=�y��ؾXeF����Cq�2�i|���M�"��z�-��&�� �.KH�)/?�:V���>6�k0?��RB���_�0Ծ�R5�����O�ӑ�&�\�3�{rny�{������F�m���Ay��7�;a,XH7~I�g>ؓG�[u"�c6�*V
�]WGm��0�sR�8ď����<#N�XG�����W;�Z]mT�M>ʴ� �L7ڂW�$ 8�L�o�9�7�gL3���I_K�g~��KI�2<'����P�}���`sf$Tt(���(	�'�S��>:��X���Y���V�̐�U32��Ee���zOmE�����؉�P'D�$ذͬ�)p%�Pj~r���+̪X��ۂ:V=K�9R:�����{;��̣֌���fE|8�tz̚�)�y��8򤄽��\<�*s!�LϹ�8k�����*k߱{%9��@)�՗���h�f����Ƚр�`��9��������W9�u�P�P�kU�4>FG4������i���<�
���`�9t�b�q%�f���I�1�j�``��=��o?j�-׏Md*����8���e�"����|!Bo��4�P4�q�}��0F>^.J�����M�ev^��ב���,��DyLϺkGݚe�@�C��赸V�p�7iyUP:Jc����*,���rAQu_
Փą��+�NX�k���� }N.�/���J����MWl�NYW��'w�����ݧa�����'ݣ\���Ϋ��Z��)��j��h��:���o�֖�<�,Ş�Y�b��X
�1�%W{�yJ�<0�t-���"W\�+��y���ɞ�^�]`�iK#ٶp�F�`N�0HMrY�=���lPP�<�A�OPUYJ
JF�n�)�Okr1:��v^��M�/:���Ox��)�76PWL�eY�VJ�_�_X[�߂���=⍚��^��V��N�wJ\�`/�7
~E��� A���ܸ��NETG��_����ŢWA�����p��A)
��A�"?�����~)H篪���,�3*b�M��X�~�^Ρ<���kǿ�:��}�4Ms�	m��)����"g�FsU���9�+���4��N��^5�Z	�bD[�3�)6�=��O��C����L�r�����̬󝵽<����=��*��NE�����T�# ����\�'��:���ƥ�5�-�ճ3�4�+�z���u�x�@z�AZ:d�A'>�9�A�}4�rv�zvOSNE�����[m�M���)��J�s�^:�L�"o��D�pq�K��j�z��I.��i@#�ӕaS�5��)��)`�rtH�o��`���ǵ*��bȚ��A+s�䏀�kpe�E5�1�De)$�ZC�?�*�a/ɖ#c���S� ��:�К�m$w�����顩�G����.��]��ϟ�Υ�<������$�N�k�^��2����l�f�l^�5��w�E�,u/���@	�4�s�C?VZg�ט�4�A�C~��%p1��F��L�R̋i�A�R<K��s�췠��U�LdY0��Z�KT�n
� �7M������A���`z�w�X���mX4ܸ���l���f6H�x,��!�q:
�%Qc_O�lی{�b��틮�����[o�#�7BOW��]}�I��,saA>p�{˲.��W=�/\5])��Gw�?�a�eĬ�|��*h��z�<z���C%��y��m����$Q���]qjlPW2d2>��&ً���Ӝ�-��{��Bv=�k���N�$�q�5L���	��1W��qR�����0�RB��=�a��e���§F������Jn�pϋ�� �eU��#Έ6���G��P��8��\���lB�7"5���tw�.�<���Z�:MݗIT�6�5�ɒ����״�h�G'�d���(�];��0C�<X��㺧t����OpʬO������ȝ�fa�B=v�öӭ~հ���l� �kϡ�_h�����LY�'����Q��u�#� �|i4�pAR�H���>�{�\��A�t��+4�f�б�M�*A�?� E��BB�v`O���Z����H��g�*�㢐�f��8nT�Cx\&�zho�F���k�	L�$dC�] u�_#����WM%=bn��2|������}�n;��q�:���|GO�\9�b����T��S^��bp,�➠Y*9�8�h�������z�<�@7��B�Td<�vb��c�0'HSg���q-��
a.��Ce���*j'�HI���𚷻Ć^��*�x��C4�(��y<O�$�`cIF��Z�-�F:��)9�N��<�Y̒~M\n52pv�EF��V���RـH����������h
.���lk~8��}ٜ�jh�~��߻~�z`�����9˶��^���W��3��w�;������J>s=s=�"f�3�������P����3�:N�y]�a]�<���-;7�y��� PK   $xX���^  �     jsons/user_defined.jsonřmO�:��
��[��o�+�Bw�	���4�-#�%��t!����F�.a�.M��Ǯ��p?��at4Z-C�ه,/��G�B���"��<�xe��M�������g�y��zuc�u���휩×����F#�`��4�>���+�#AFLP@V(Y���9M@O���*lB�����E���ڇ���\g�q�-�
#˽CVY���8>Y_�s��8)�rtt?*V7�|����7�<�qd�������yy���'���Ȫȿ�bŉ���<���5�e�Dz����'
�cI�Ds`:6ɗ��]�U|�i�scC�~�0ގ�4Z�Й�/��I���M�l��l�f���O������6���{���r�:_/�f!��h���k�b^���x�8����͕7��E}�$���%�+�5�r��?矝q�a=ПM�V~����)����*cXuU��jt�I�Ǒ�Ė�@l����t�QĵǐŘV���i�y,1J!f�G�B��iM�8�W�L;�#�:*ځ�2QnUPN$��k��qQ�~��o���pp��	���6Ç�i~�����__pqç����ظ����C�p��CO8M�E�{�Y.�pݓ͓l�d��l�d�$[�d˴HiQS����4<�i_Ku�v����8�$=mhOAg ���/N�]�5�k)��ӓ���.���_���\����]_��D�+�AWY��D]q��T̯����bh.���%[��C��4�xȖ���|<M�L�e�;0#O�ٞl������l������;��𶧶SH�wX�S�i:s���Tvz~�6��alOa�Վ/v����2=�x�wz�׵�m������L��wǟ?~Hw����cѯ��u�u�k;�����O�u��q71��n_Y�z�&2t�͋xk�=���O��eQ<6���Eє��|�>C7a�&�8���D{]޾/���&���|�/s;�kU��Zw�>'6����̸zUœ�]�'�=t�S�8/��q�1))�(��1L���A諃?M]���E�Cy���C�1K="�Sd�1HJʑ�$7A2�����Xz'�bJ�A[�q�R,$�4��q��3�c�0@�2��bY�%r$�Fd܂�}��tB((�V� 0����uXq"n����,b��=��@�'~����z{�K�?�)^ ��ɪU^�~�<�ދ�{����-a�0D��Uϵ֊g�#'l�X&�ye��Lp&d��ז�3�͚J!�M�/j���X!�ɤ7�uT��1��Yh�VQ��4	! ��C;�l��b� Tl��$*�_�!!zBPGK����b?Ez�K���lo�-e�����6l�]xw���X�����
y��?/>=|PK
   $xXkU���  ��                  cirkitFile.jsonPK
   $xXo�>��q  �q  /             !  images/2cd737db-51bc-41eb-8762-f3273c40eae5.pngPK
   �zxX;��d  �)  /             8�  images/35440911-0bff-4ebf-83cc-bd2192eee111.pngPK
   $xX����+  J  /             �  images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.pngPK
   ��WǆO2K 9X /             a�  images/59f150f1-5697-4080-b5dc-b8b306a70e65.pngPK
   ��WǆO2K 9X /             �� images/83b09b1d-e584-4d9e-8c7e-ad4061c788ce.pngPK
   $xXN�v4	� m� /             %K images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.pngPK
   $xX~��a� ٮ /             { images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.pngPK
   �zxXp+��  y4  /             )� images/f9f29454-e4d8-4baa-8657-cb66eaf7dadc.pngPK
   $xX���^  �               b� jsons/user_defined.jsonPK    
 
 j  ��   